------------------------------------------------------------
-- VHDL TK510_Mekanisk
-- 2017 1 13 17 4 7
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.0.6.282
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK510_Mekanisk
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK510_Mekanisk Is
  attribute MacroCell : boolean;

End TK510_Mekanisk;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK510_Mekanisk Is
   Component X_2392                                          -- ObjectKind=Part|PrimaryId=M51000|SecondaryId=1
   End Component;



   attribute antall : string;
   attribute antall of M51017 : Label is "30";
   attribute antall of M51016 : Label is "30";
   attribute antall of M51015 : Label is "30";
   attribute antall of M51014 : Label is "30";
   attribute antall of M51013 : Label is "30";
   attribute antall of M51012 : Label is "30";
   attribute antall of M51011 : Label is "30";
   attribute antall of M51010 : Label is "30";
   attribute antall of M51009 : Label is "30";
   attribute antall of M51008 : Label is "30";
   attribute antall of M51007 : Label is "30";
   attribute antall of M51006 : Label is "30";
   attribute antall of M51005 : Label is "30";
   attribute antall of M51004 : Label is "30";
   attribute antall of M51003 : Label is "30";
   attribute antall of M51002 : Label is "30";
   attribute antall of M51001 : Label is "30";
   attribute antall of M51000 : Label is "30";

   attribute Database_Table_Name : string;
   attribute Database_Table_Name of M51017 : Label is "altium";
   attribute Database_Table_Name of M51016 : Label is "altium";
   attribute Database_Table_Name of M51015 : Label is "altium";
   attribute Database_Table_Name of M51014 : Label is "altium";
   attribute Database_Table_Name of M51013 : Label is "altium";
   attribute Database_Table_Name of M51012 : Label is "altium";
   attribute Database_Table_Name of M51011 : Label is "altium";
   attribute Database_Table_Name of M51010 : Label is "altium";
   attribute Database_Table_Name of M51009 : Label is "altium";
   attribute Database_Table_Name of M51008 : Label is "altium";
   attribute Database_Table_Name of M51007 : Label is "altium";
   attribute Database_Table_Name of M51006 : Label is "altium";
   attribute Database_Table_Name of M51005 : Label is "altium";
   attribute Database_Table_Name of M51004 : Label is "altium";
   attribute Database_Table_Name of M51003 : Label is "altium";
   attribute Database_Table_Name of M51002 : Label is "altium";
   attribute Database_Table_Name of M51001 : Label is "altium";
   attribute Database_Table_Name of M51000 : Label is "altium";

   attribute dybde : string;
   attribute dybde of M51017 : Label is "0";
   attribute dybde of M51016 : Label is "0";
   attribute dybde of M51015 : Label is "0";
   attribute dybde of M51014 : Label is "0";
   attribute dybde of M51013 : Label is "0";
   attribute dybde of M51012 : Label is "0";
   attribute dybde of M51011 : Label is "0";
   attribute dybde of M51010 : Label is "0";
   attribute dybde of M51009 : Label is "0";
   attribute dybde of M51008 : Label is "0";
   attribute dybde of M51007 : Label is "0";
   attribute dybde of M51006 : Label is "0";
   attribute dybde of M51005 : Label is "0";
   attribute dybde of M51004 : Label is "0";
   attribute dybde of M51003 : Label is "0";
   attribute dybde of M51002 : Label is "0";
   attribute dybde of M51001 : Label is "0";
   attribute dybde of M51000 : Label is "0";

   attribute hylle : string;
   attribute hylle of M51017 : Label is "15";
   attribute hylle of M51016 : Label is "15";
   attribute hylle of M51015 : Label is "15";
   attribute hylle of M51014 : Label is "15";
   attribute hylle of M51013 : Label is "15";
   attribute hylle of M51012 : Label is "15";
   attribute hylle of M51011 : Label is "15";
   attribute hylle of M51010 : Label is "15";
   attribute hylle of M51009 : Label is "15";
   attribute hylle of M51008 : Label is "15";
   attribute hylle of M51007 : Label is "15";
   attribute hylle of M51006 : Label is "15";
   attribute hylle of M51005 : Label is "15";
   attribute hylle of M51004 : Label is "15";
   attribute hylle of M51003 : Label is "15";
   attribute hylle of M51002 : Label is "15";
   attribute hylle of M51001 : Label is "15";
   attribute hylle of M51000 : Label is "15";

   attribute id : string;
   attribute id of M51017 : Label is "2392";
   attribute id of M51016 : Label is "2392";
   attribute id of M51015 : Label is "2392";
   attribute id of M51014 : Label is "2392";
   attribute id of M51013 : Label is "2392";
   attribute id of M51012 : Label is "2392";
   attribute id of M51011 : Label is "2392";
   attribute id of M51010 : Label is "2392";
   attribute id of M51009 : Label is "2392";
   attribute id of M51008 : Label is "2392";
   attribute id of M51007 : Label is "2392";
   attribute id of M51006 : Label is "2392";
   attribute id of M51005 : Label is "2392";
   attribute id of M51004 : Label is "2392";
   attribute id of M51003 : Label is "2392";
   attribute id of M51002 : Label is "2392";
   attribute id of M51001 : Label is "2392";
   attribute id of M51000 : Label is "2392";

   attribute kolonne : string;
   attribute kolonne of M51017 : Label is "2";
   attribute kolonne of M51016 : Label is "2";
   attribute kolonne of M51015 : Label is "2";
   attribute kolonne of M51014 : Label is "2";
   attribute kolonne of M51013 : Label is "2";
   attribute kolonne of M51012 : Label is "2";
   attribute kolonne of M51011 : Label is "2";
   attribute kolonne of M51010 : Label is "2";
   attribute kolonne of M51009 : Label is "2";
   attribute kolonne of M51008 : Label is "2";
   attribute kolonne of M51007 : Label is "2";
   attribute kolonne of M51006 : Label is "2";
   attribute kolonne of M51005 : Label is "2";
   attribute kolonne of M51004 : Label is "2";
   attribute kolonne of M51003 : Label is "2";
   attribute kolonne of M51002 : Label is "2";
   attribute kolonne of M51001 : Label is "2";
   attribute kolonne of M51000 : Label is "2";

   attribute lager_type : string;
   attribute lager_type of M51017 : Label is "Fremlager";
   attribute lager_type of M51016 : Label is "Fremlager";
   attribute lager_type of M51015 : Label is "Fremlager";
   attribute lager_type of M51014 : Label is "Fremlager";
   attribute lager_type of M51013 : Label is "Fremlager";
   attribute lager_type of M51012 : Label is "Fremlager";
   attribute lager_type of M51011 : Label is "Fremlager";
   attribute lager_type of M51010 : Label is "Fremlager";
   attribute lager_type of M51009 : Label is "Fremlager";
   attribute lager_type of M51008 : Label is "Fremlager";
   attribute lager_type of M51007 : Label is "Fremlager";
   attribute lager_type of M51006 : Label is "Fremlager";
   attribute lager_type of M51005 : Label is "Fremlager";
   attribute lager_type of M51004 : Label is "Fremlager";
   attribute lager_type of M51003 : Label is "Fremlager";
   attribute lager_type of M51002 : Label is "Fremlager";
   attribute lager_type of M51001 : Label is "Fremlager";
   attribute lager_type of M51000 : Label is "Fremlager";

   attribute navn : string;
   attribute navn of M51017 : Label is "KortSt�tte";
   attribute navn of M51016 : Label is "KortSt�tte";
   attribute navn of M51015 : Label is "KortSt�tte";
   attribute navn of M51014 : Label is "KortSt�tte";
   attribute navn of M51013 : Label is "KortSt�tte";
   attribute navn of M51012 : Label is "KortSt�tte";
   attribute navn of M51011 : Label is "KortSt�tte";
   attribute navn of M51010 : Label is "KortSt�tte";
   attribute navn of M51009 : Label is "KortSt�tte";
   attribute navn of M51008 : Label is "KortSt�tte";
   attribute navn of M51007 : Label is "KortSt�tte";
   attribute navn of M51006 : Label is "KortSt�tte";
   attribute navn of M51005 : Label is "KortSt�tte";
   attribute navn of M51004 : Label is "KortSt�tte";
   attribute navn of M51003 : Label is "KortSt�tte";
   attribute navn of M51002 : Label is "KortSt�tte";
   attribute navn of M51001 : Label is "KortSt�tte";
   attribute navn of M51000 : Label is "KortSt�tte";

   attribute nokkelord : string;
   attribute nokkelord of M51017 : Label is "support";
   attribute nokkelord of M51016 : Label is "support";
   attribute nokkelord of M51015 : Label is "support";
   attribute nokkelord of M51014 : Label is "support";
   attribute nokkelord of M51013 : Label is "support";
   attribute nokkelord of M51012 : Label is "support";
   attribute nokkelord of M51011 : Label is "support";
   attribute nokkelord of M51010 : Label is "support";
   attribute nokkelord of M51009 : Label is "support";
   attribute nokkelord of M51008 : Label is "support";
   attribute nokkelord of M51007 : Label is "support";
   attribute nokkelord of M51006 : Label is "support";
   attribute nokkelord of M51005 : Label is "support";
   attribute nokkelord of M51004 : Label is "support";
   attribute nokkelord of M51003 : Label is "support";
   attribute nokkelord of M51002 : Label is "support";
   attribute nokkelord of M51001 : Label is "support";
   attribute nokkelord of M51000 : Label is "support";

   attribute pakke_opprettet : string;
   attribute pakke_opprettet of M51017 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51016 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51015 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51014 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51013 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51012 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51011 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51010 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51009 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51008 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51007 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51006 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51005 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51004 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51003 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51002 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51001 : Label is "12.07.2014 20.29.43";
   attribute pakke_opprettet of M51000 : Label is "12.07.2014 20.29.43";

   attribute pakke_opprettet_av : string;
   attribute pakke_opprettet_av of M51017 : Label is "815";
   attribute pakke_opprettet_av of M51016 : Label is "815";
   attribute pakke_opprettet_av of M51015 : Label is "815";
   attribute pakke_opprettet_av of M51014 : Label is "815";
   attribute pakke_opprettet_av of M51013 : Label is "815";
   attribute pakke_opprettet_av of M51012 : Label is "815";
   attribute pakke_opprettet_av of M51011 : Label is "815";
   attribute pakke_opprettet_av of M51010 : Label is "815";
   attribute pakke_opprettet_av of M51009 : Label is "815";
   attribute pakke_opprettet_av of M51008 : Label is "815";
   attribute pakke_opprettet_av of M51007 : Label is "815";
   attribute pakke_opprettet_av of M51006 : Label is "815";
   attribute pakke_opprettet_av of M51005 : Label is "815";
   attribute pakke_opprettet_av of M51004 : Label is "815";
   attribute pakke_opprettet_av of M51003 : Label is "815";
   attribute pakke_opprettet_av of M51002 : Label is "815";
   attribute pakke_opprettet_av of M51001 : Label is "815";
   attribute pakke_opprettet_av of M51000 : Label is "815";

   attribute pakketype : string;
   attribute pakketype of M51017 : Label is "TH";
   attribute pakketype of M51016 : Label is "TH";
   attribute pakketype of M51015 : Label is "TH";
   attribute pakketype of M51014 : Label is "TH";
   attribute pakketype of M51013 : Label is "TH";
   attribute pakketype of M51012 : Label is "TH";
   attribute pakketype of M51011 : Label is "TH";
   attribute pakketype of M51010 : Label is "TH";
   attribute pakketype of M51009 : Label is "TH";
   attribute pakketype of M51008 : Label is "TH";
   attribute pakketype of M51007 : Label is "TH";
   attribute pakketype of M51006 : Label is "TH";
   attribute pakketype of M51005 : Label is "TH";
   attribute pakketype of M51004 : Label is "TH";
   attribute pakketype of M51003 : Label is "TH";
   attribute pakketype of M51002 : Label is "TH";
   attribute pakketype of M51001 : Label is "TH";
   attribute pakketype of M51000 : Label is "TH";

   attribute pris : string;
   attribute pris of M51017 : Label is "5";
   attribute pris of M51016 : Label is "5";
   attribute pris of M51015 : Label is "5";
   attribute pris of M51014 : Label is "5";
   attribute pris of M51013 : Label is "5";
   attribute pris of M51012 : Label is "5";
   attribute pris of M51011 : Label is "5";
   attribute pris of M51010 : Label is "5";
   attribute pris of M51009 : Label is "5";
   attribute pris of M51008 : Label is "5";
   attribute pris of M51007 : Label is "5";
   attribute pris of M51006 : Label is "5";
   attribute pris of M51005 : Label is "5";
   attribute pris of M51004 : Label is "5";
   attribute pris of M51003 : Label is "5";
   attribute pris of M51002 : Label is "5";
   attribute pris of M51001 : Label is "5";
   attribute pris of M51000 : Label is "5";

   attribute rad : string;
   attribute rad of M51017 : Label is "5";
   attribute rad of M51016 : Label is "5";
   attribute rad of M51015 : Label is "5";
   attribute rad of M51014 : Label is "5";
   attribute rad of M51013 : Label is "5";
   attribute rad of M51012 : Label is "5";
   attribute rad of M51011 : Label is "5";
   attribute rad of M51010 : Label is "5";
   attribute rad of M51009 : Label is "5";
   attribute rad of M51008 : Label is "5";
   attribute rad of M51007 : Label is "5";
   attribute rad of M51006 : Label is "5";
   attribute rad of M51005 : Label is "5";
   attribute rad of M51004 : Label is "5";
   attribute rad of M51003 : Label is "5";
   attribute rad of M51002 : Label is "5";
   attribute rad of M51001 : Label is "5";
   attribute rad of M51000 : Label is "5";

   attribute rom : string;
   attribute rom of M51017 : Label is "OV";
   attribute rom of M51016 : Label is "OV";
   attribute rom of M51015 : Label is "OV";
   attribute rom of M51014 : Label is "OV";
   attribute rom of M51013 : Label is "OV";
   attribute rom of M51012 : Label is "OV";
   attribute rom of M51011 : Label is "OV";
   attribute rom of M51010 : Label is "OV";
   attribute rom of M51009 : Label is "OV";
   attribute rom of M51008 : Label is "OV";
   attribute rom of M51007 : Label is "OV";
   attribute rom of M51006 : Label is "OV";
   attribute rom of M51005 : Label is "OV";
   attribute rom of M51004 : Label is "OV";
   attribute rom of M51003 : Label is "OV";
   attribute rom of M51002 : Label is "OV";
   attribute rom of M51001 : Label is "OV";
   attribute rom of M51000 : Label is "OV";

   attribute symbol_opprettet : string;
   attribute symbol_opprettet of M51017 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51016 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51015 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51014 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51013 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51012 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51011 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51010 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51009 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51008 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51007 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51006 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51005 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51004 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51003 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51002 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51001 : Label is "12.07.2014 20.29.53";
   attribute symbol_opprettet of M51000 : Label is "12.07.2014 20.29.53";

   attribute symbol_opprettet_av : string;
   attribute symbol_opprettet_av of M51017 : Label is "815";
   attribute symbol_opprettet_av of M51016 : Label is "815";
   attribute symbol_opprettet_av of M51015 : Label is "815";
   attribute symbol_opprettet_av of M51014 : Label is "815";
   attribute symbol_opprettet_av of M51013 : Label is "815";
   attribute symbol_opprettet_av of M51012 : Label is "815";
   attribute symbol_opprettet_av of M51011 : Label is "815";
   attribute symbol_opprettet_av of M51010 : Label is "815";
   attribute symbol_opprettet_av of M51009 : Label is "815";
   attribute symbol_opprettet_av of M51008 : Label is "815";
   attribute symbol_opprettet_av of M51007 : Label is "815";
   attribute symbol_opprettet_av of M51006 : Label is "815";
   attribute symbol_opprettet_av of M51005 : Label is "815";
   attribute symbol_opprettet_av of M51004 : Label is "815";
   attribute symbol_opprettet_av of M51003 : Label is "815";
   attribute symbol_opprettet_av of M51002 : Label is "815";
   attribute symbol_opprettet_av of M51001 : Label is "815";
   attribute symbol_opprettet_av of M51000 : Label is "815";


Begin
    M51017 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51017|SecondaryId=1
;

    M51016 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51016|SecondaryId=1
;

    M51015 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51015|SecondaryId=1
;

    M51014 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51014|SecondaryId=1
;

    M51013 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51013|SecondaryId=1
;

    M51012 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51012|SecondaryId=1
;

    M51011 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51011|SecondaryId=1
;

    M51010 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51010|SecondaryId=1
;

    M51009 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51009|SecondaryId=1
;

    M51008 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51008|SecondaryId=1
;

    M51007 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51007|SecondaryId=1
;

    M51006 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51006|SecondaryId=1
;

    M51005 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51005|SecondaryId=1
;

    M51004 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51004|SecondaryId=1
;

    M51003 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51003|SecondaryId=1
;

    M51002 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51002|SecondaryId=1
;

    M51001 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51001|SecondaryId=1
;

    M51000 : X_2392                                          -- ObjectKind=Part|PrimaryId=M51000|SecondaryId=1
;

End Structure;
------------------------------------------------------------

