------------------------------------------------------------
-- VHDL TK510_Kontakter
-- 2014 7 6 17 49 11
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.11.33708
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK510_Kontakter
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK510_Kontakter Is
  attribute MacroCell : boolean;

End TK510_Kontakter;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK510_Kontakter Is
   Component PCI_ExpressMINUS36P                             -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
      port
      (
        A1  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A1
        A2  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A2
        A3  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A3
        A4  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A4
        A5  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A5
        A6  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A6
        A7  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A7
        A8  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A8
        A9  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A9
        A10 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A10
        A11 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A11
        A12 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A12
        A13 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A13
        A14 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A14
        A15 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A15
        A16 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A16
        A17 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A17
        A18 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-A18
        B1  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B1
        B2  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B2
        B3  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B3
        B4  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B4
        B5  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B5
        B6  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B6
        B7  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B7
        B8  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B8
        B9  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B9
        B10 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B10
        B11 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B11
        B12 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B12
        B13 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B13
        B14 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B14
        B15 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B15
        B16 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B16
        B17 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J?-B17
        B18 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=J?-B18
      );
   End Component;



   attribute beskrivelse : string;
   attribute beskrivelse of J? : Label is "PCI_Express-36P";

   attribute Database_Table_Name : string;
   attribute Database_Table_Name of J? : Label is "altium";

   attribute leverandor : string;
   attribute leverandor of J? : Label is "Farnell";

   attribute leverandor_varenr : string;
   attribute leverandor_varenr of J? : Label is "1144435";

   attribute navn : string;
   attribute navn of J? : Label is "PCI_Express-36P";

   attribute nokkelord : string;
   attribute nokkelord of J? : Label is "Card-edge";

   attribute pakke_opprettet : string;
   attribute pakke_opprettet of J? : Label is "06.07.2014 17:26:47";

   attribute pakke_opprettet_av : string;
   attribute pakke_opprettet_av of J? : Label is "815";

   attribute pakketype : string;
   attribute pakketype of J? : Label is "92";

   attribute pris : string;
   attribute pris of J? : Label is "16";

   attribute produsent : string;
   attribute produsent of J? : Label is "FCI";

   attribute symbol_opprettet : string;
   attribute symbol_opprettet of J? : Label is "06.07.2014 17:26:37";

   attribute symbol_opprettet_av : string;
   attribute symbol_opprettet_av of J? : Label is "815";


Begin
    J : PCI_ExpressMINUS36P                                  -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
;

    J : PCI_ExpressMINUS36P                                  -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
;

    J : PCI_ExpressMINUS36P                                  -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
;

    J : PCI_ExpressMINUS36P                                  -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
;

    J : PCI_ExpressMINUS36P                                  -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
;

    J : PCI_ExpressMINUS36P                                  -- ObjectKind=Part|PrimaryId=J?|SecondaryId=1
;

End Structure;
------------------------------------------------------------

