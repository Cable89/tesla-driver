------------------------------------------------------------
-- VHDL TK510_Spenningsforsyninger
-- 2017 1 13 17 4 10
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.0.6.282
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK510_Spenningsforsyninger
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK510_Spenningsforsyninger Is
  port
  (
    BUS_B5           : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B5
    BUS_B6           : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B6
    BUS_B7           : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B7
    BUS_B8           : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B8
    BUS_B9           : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B9
    BUS_B10          : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B10
    BUS_B11          : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.B11
    BUS_INTERRUPT    : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.INTERRUPT
    BUS_KORT_INNSATT : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.KORT_INNSATT
    BUS_LIMIT        : InOut STD_LOGIC;                      -- ObjectKind=Port|PrimaryId=BUS.LIMIT
    BUS_TRIGGER      : InOut STD_LOGIC                       -- ObjectKind=Port|PrimaryId=BUS.TRIGGER
  );
  attribute MacroCell : boolean;

End TK510_Spenningsforsyninger;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK510_Spenningsforsyninger Is
   Component X_2209                                          -- ObjectKind=Part|PrimaryId=D51001|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=D51001-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=D51001-2
      );
   End Component;

   Component X_2212                                          -- ObjectKind=Part|PrimaryId=Q51016|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=Q51016-1
        X_2 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=Q51016-2
        X_3 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=Q51016-3
      );
   End Component;

   Component X_2213                                          -- ObjectKind=Part|PrimaryId=Q51013|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=Q51013-1
        X_2 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=Q51013-2
        X_3 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=Q51013-3
      );
   End Component;

   Component X_2227                                          -- ObjectKind=Part|PrimaryId=J51029|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51029-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=J51029-2
      );
   End Component;

   Component X_2382                                          -- ObjectKind=Part|PrimaryId=J51007|SecondaryId=1
      port
      (
        A1  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A1
        A2  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A2
        A3  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A3
        A4  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A4
        A5  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A5
        A6  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A6
        A7  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A7
        A8  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A8
        A9  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A9
        A10 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A10
        A11 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A11
        A12 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A12
        A13 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A13
        A14 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A14
        A15 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A15
        A16 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A16
        A17 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A17
        A18 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-A18
        B1  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B1
        B2  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B2
        B3  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B3
        B4  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B4
        B5  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B5
        B6  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B6
        B7  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B7
        B8  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B8
        B9  : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B9
        B10 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B10
        B11 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B11
        B12 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B12
        B13 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B13
        B14 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B14
        B15 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B15
        B16 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B16
        B17 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J51007-B17
        B18 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=J51007-B18
      );
   End Component;

   Component X_2444                                          -- ObjectKind=Part|PrimaryId=R51041|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=R51041-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=R51041-2
      );
   End Component;

   Component X_2448                                          -- ObjectKind=Part|PrimaryId=R51044|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=R51044-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=R51044-2
      );
   End Component;


    Signal NamedSignal_AC_S6_L1        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=AC_S6_L1
    Signal NamedSignal_AC_S6_L2        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=AC_S6_L2
    Signal NamedSignal_AC_S7_L1        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=AC_S7_L1
    Signal NamedSignal_AC_S7_L2        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=AC_S7_L2
    Signal NamedSignal_AC_S8_L1        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=AC_S8_L1
    Signal NamedSignal_AC_S8_L2        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=AC_S8_L2
    Signal PinSignal_D51001_1          : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD51001_1
    Signal PinSignal_D51002_1          : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD51002_1
    Signal PinSignal_D51003_1          : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD51003_1
    Signal PinSignal_J51007_A1         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    Signal PinSignal_J51007_A10        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    Signal PinSignal_J51007_A11        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    Signal PinSignal_J51007_A2         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    Signal PinSignal_J51007_A3         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    Signal PinSignal_J51007_A4         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    Signal PinSignal_J51007_A5         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    Signal PinSignal_J51007_A6         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    Signal PinSignal_J51007_A7         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    Signal PinSignal_J51007_A8         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    Signal PinSignal_J51007_A9         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    Signal PinSignal_J51007_B1         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51007_B1
    Signal PinSignal_J51008_A1         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    Signal PinSignal_J51008_A10        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    Signal PinSignal_J51008_A11        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    Signal PinSignal_J51008_A2         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    Signal PinSignal_J51008_A3         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    Signal PinSignal_J51008_A4         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    Signal PinSignal_J51008_A5         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    Signal PinSignal_J51008_A6         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    Signal PinSignal_J51008_A7         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    Signal PinSignal_J51008_A8         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    Signal PinSignal_J51008_A9         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    Signal PinSignal_J51008_B1         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51008_B1
    Signal PinSignal_J51028_A1         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    Signal PinSignal_J51028_A10        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    Signal PinSignal_J51028_A11        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    Signal PinSignal_J51028_A2         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    Signal PinSignal_J51028_A3         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    Signal PinSignal_J51028_A4         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    Signal PinSignal_J51028_A5         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    Signal PinSignal_J51028_A6         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    Signal PinSignal_J51028_A7         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    Signal PinSignal_J51028_A8         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    Signal PinSignal_J51028_A9         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    Signal PinSignal_J51028_B1         : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ51028_B1
    Signal PinSignal_Q51016_2          : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetQ51016_2
    Signal PinSignal_Q51017_2          : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetQ51017_2
    Signal PinSignal_Q51018_2          : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetQ51018_2
    Signal PowerSignal_GND             : STD_LOGIC; -- ObjectKind=Net|PrimaryId=GND
    Signal PowerSignal_VCC_EXTRA       : STD_LOGIC; -- ObjectKind=Net|PrimaryId=VCC_EXTRA
    Signal PowerSignal_VCC_P18V        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=VCC_P18V
    Signal PowerSignal_VCC_P5V0        : STD_LOGIC; -- ObjectKind=Net|PrimaryId=VCC_P5V0

   attribute antall : string;
   attribute antall of R51046 : Label is "100";
   attribute antall of R51045 : Label is "100";
   attribute antall of R51044 : Label is "100";
   attribute antall of R51043 : Label is "100";
   attribute antall of R51042 : Label is "100";
   attribute antall of R51041 : Label is "100";
   attribute antall of Q51015 : Label is "100";
   attribute antall of Q51014 : Label is "100";
   attribute antall of Q51013 : Label is "100";
   attribute antall of J51049 : Label is "100";
   attribute antall of J51048 : Label is "100";
   attribute antall of J51047 : Label is "100";
   attribute antall of J51046 : Label is "100";
   attribute antall of J51045 : Label is "100";
   attribute antall of J51044 : Label is "100";
   attribute antall of J51043 : Label is "100";
   attribute antall of J51042 : Label is "100";
   attribute antall of J51041 : Label is "100";
   attribute antall of J51040 : Label is "100";
   attribute antall of J51039 : Label is "100";
   attribute antall of J51038 : Label is "100";
   attribute antall of J51037 : Label is "100";
   attribute antall of J51036 : Label is "100";
   attribute antall of J51035 : Label is "100";
   attribute antall of J51034 : Label is "100";
   attribute antall of J51033 : Label is "100";
   attribute antall of J51032 : Label is "100";
   attribute antall of J51031 : Label is "100";
   attribute antall of J51030 : Label is "100";
   attribute antall of J51029 : Label is "100";
   attribute antall of D51003 : Label is "50";
   attribute antall of D51002 : Label is "50";
   attribute antall of D51001 : Label is "50";

   attribute beskrivelse : string;
   attribute beskrivelse of D51003 : Label is "SMD";
   attribute beskrivelse of D51002 : Label is "SMD";
   attribute beskrivelse of D51001 : Label is "SMD";

   attribute Database_Table_Name : string;
   attribute Database_Table_Name of R51046 : Label is "altium_Motstander";
   attribute Database_Table_Name of R51045 : Label is "altium_Motstander";
   attribute Database_Table_Name of R51044 : Label is "altium_Motstander";
   attribute Database_Table_Name of R51043 : Label is "altium_Motstander";
   attribute Database_Table_Name of R51042 : Label is "altium_Motstander";
   attribute Database_Table_Name of R51041 : Label is "altium_Motstander";
   attribute Database_Table_Name of Q51018 : Label is "altium_Transistorer";
   attribute Database_Table_Name of Q51017 : Label is "altium_Transistorer";
   attribute Database_Table_Name of Q51016 : Label is "altium_Transistorer";
   attribute Database_Table_Name of Q51015 : Label is "altium_Transistorer";
   attribute Database_Table_Name of Q51014 : Label is "altium_Transistorer";
   attribute Database_Table_Name of Q51013 : Label is "altium_Transistorer";
   attribute Database_Table_Name of J51049 : Label is "altium";
   attribute Database_Table_Name of J51048 : Label is "altium";
   attribute Database_Table_Name of J51047 : Label is "altium";
   attribute Database_Table_Name of J51046 : Label is "altium";
   attribute Database_Table_Name of J51045 : Label is "altium";
   attribute Database_Table_Name of J51044 : Label is "altium";
   attribute Database_Table_Name of J51043 : Label is "altium";
   attribute Database_Table_Name of J51042 : Label is "altium";
   attribute Database_Table_Name of J51041 : Label is "altium";
   attribute Database_Table_Name of J51040 : Label is "altium";
   attribute Database_Table_Name of J51039 : Label is "altium";
   attribute Database_Table_Name of J51038 : Label is "altium";
   attribute Database_Table_Name of J51037 : Label is "altium";
   attribute Database_Table_Name of J51036 : Label is "altium";
   attribute Database_Table_Name of J51035 : Label is "altium";
   attribute Database_Table_Name of J51034 : Label is "altium";
   attribute Database_Table_Name of J51033 : Label is "altium";
   attribute Database_Table_Name of J51032 : Label is "altium";
   attribute Database_Table_Name of J51031 : Label is "altium";
   attribute Database_Table_Name of J51030 : Label is "altium";
   attribute Database_Table_Name of J51029 : Label is "altium";
   attribute Database_Table_Name of J51028 : Label is "altium";
   attribute Database_Table_Name of J51008 : Label is "altium";
   attribute Database_Table_Name of J51007 : Label is "altium";
   attribute Database_Table_Name of D51003 : Label is "altium_Dioder";
   attribute Database_Table_Name of D51002 : Label is "altium_Dioder";
   attribute Database_Table_Name of D51001 : Label is "altium_Dioder";

   attribute Design_comment : string;
   attribute Design_comment of Q51018 : Label is "";
   attribute Design_comment of Q51017 : Label is "";
   attribute Design_comment of Q51016 : Label is "";

   attribute dybde : string;
   attribute dybde of R51046 : Label is "36";
   attribute dybde of R51045 : Label is "36";
   attribute dybde of R51044 : Label is "36";
   attribute dybde of R51043 : Label is "72";
   attribute dybde of R51042 : Label is "72";
   attribute dybde of R51041 : Label is "72";
   attribute dybde of Q51015 : Label is "0";
   attribute dybde of Q51014 : Label is "0";
   attribute dybde of Q51013 : Label is "0";
   attribute dybde of J51049 : Label is "0";
   attribute dybde of J51048 : Label is "0";
   attribute dybde of J51047 : Label is "0";
   attribute dybde of J51046 : Label is "0";
   attribute dybde of J51045 : Label is "0";
   attribute dybde of J51044 : Label is "0";
   attribute dybde of J51043 : Label is "0";
   attribute dybde of J51042 : Label is "0";
   attribute dybde of J51041 : Label is "0";
   attribute dybde of J51040 : Label is "0";
   attribute dybde of J51039 : Label is "0";
   attribute dybde of J51038 : Label is "0";
   attribute dybde of J51037 : Label is "0";
   attribute dybde of J51036 : Label is "0";
   attribute dybde of J51035 : Label is "0";
   attribute dybde of J51034 : Label is "0";
   attribute dybde of J51033 : Label is "0";
   attribute dybde of J51032 : Label is "0";
   attribute dybde of J51031 : Label is "0";
   attribute dybde of J51030 : Label is "0";
   attribute dybde of J51029 : Label is "0";
   attribute dybde of D51003 : Label is "2";
   attribute dybde of D51002 : Label is "2";
   attribute dybde of D51001 : Label is "2";

   attribute hylle : string;
   attribute hylle of R51046 : Label is "6";
   attribute hylle of R51045 : Label is "6";
   attribute hylle of R51044 : Label is "6";
   attribute hylle of R51043 : Label is "6";
   attribute hylle of R51042 : Label is "6";
   attribute hylle of R51041 : Label is "6";
   attribute hylle of Q51015 : Label is "4";
   attribute hylle of Q51014 : Label is "4";
   attribute hylle of Q51013 : Label is "4";
   attribute hylle of J51049 : Label is "10";
   attribute hylle of J51048 : Label is "10";
   attribute hylle of J51047 : Label is "10";
   attribute hylle of J51046 : Label is "10";
   attribute hylle of J51045 : Label is "10";
   attribute hylle of J51044 : Label is "10";
   attribute hylle of J51043 : Label is "10";
   attribute hylle of J51042 : Label is "10";
   attribute hylle of J51041 : Label is "10";
   attribute hylle of J51040 : Label is "10";
   attribute hylle of J51039 : Label is "10";
   attribute hylle of J51038 : Label is "10";
   attribute hylle of J51037 : Label is "10";
   attribute hylle of J51036 : Label is "10";
   attribute hylle of J51035 : Label is "10";
   attribute hylle of J51034 : Label is "10";
   attribute hylle of J51033 : Label is "10";
   attribute hylle of J51032 : Label is "10";
   attribute hylle of J51031 : Label is "10";
   attribute hylle of J51030 : Label is "10";
   attribute hylle of J51029 : Label is "10";
   attribute hylle of D51003 : Label is "13";
   attribute hylle of D51002 : Label is "13";
   attribute hylle of D51001 : Label is "13";

   attribute id : string;
   attribute id of R51046 : Label is "2448";
   attribute id of R51045 : Label is "2448";
   attribute id of R51044 : Label is "2448";
   attribute id of R51043 : Label is "2444";
   attribute id of R51042 : Label is "2444";
   attribute id of R51041 : Label is "2444";
   attribute id of Q51018 : Label is "2212";
   attribute id of Q51017 : Label is "2212";
   attribute id of Q51016 : Label is "2212";
   attribute id of Q51015 : Label is "2213";
   attribute id of Q51014 : Label is "2213";
   attribute id of Q51013 : Label is "2213";
   attribute id of J51049 : Label is "2227";
   attribute id of J51048 : Label is "2227";
   attribute id of J51047 : Label is "2227";
   attribute id of J51046 : Label is "2227";
   attribute id of J51045 : Label is "2227";
   attribute id of J51044 : Label is "2227";
   attribute id of J51043 : Label is "2227";
   attribute id of J51042 : Label is "2227";
   attribute id of J51041 : Label is "2227";
   attribute id of J51040 : Label is "2227";
   attribute id of J51039 : Label is "2227";
   attribute id of J51038 : Label is "2227";
   attribute id of J51037 : Label is "2227";
   attribute id of J51036 : Label is "2227";
   attribute id of J51035 : Label is "2227";
   attribute id of J51034 : Label is "2227";
   attribute id of J51033 : Label is "2227";
   attribute id of J51032 : Label is "2227";
   attribute id of J51031 : Label is "2227";
   attribute id of J51030 : Label is "2227";
   attribute id of J51029 : Label is "2227";
   attribute id of J51028 : Label is "2382";
   attribute id of J51008 : Label is "2382";
   attribute id of J51007 : Label is "2382";
   attribute id of D51003 : Label is "2209";
   attribute id of D51002 : Label is "2209";
   attribute id of D51001 : Label is "2209";

   attribute kolonne : string;
   attribute kolonne of R51046 : Label is "0";
   attribute kolonne of R51045 : Label is "0";
   attribute kolonne of R51044 : Label is "0";
   attribute kolonne of R51043 : Label is "0";
   attribute kolonne of R51042 : Label is "0";
   attribute kolonne of R51041 : Label is "0";
   attribute kolonne of Q51015 : Label is "3";
   attribute kolonne of Q51014 : Label is "3";
   attribute kolonne of Q51013 : Label is "3";
   attribute kolonne of J51049 : Label is "0";
   attribute kolonne of J51048 : Label is "0";
   attribute kolonne of J51047 : Label is "0";
   attribute kolonne of J51046 : Label is "0";
   attribute kolonne of J51045 : Label is "0";
   attribute kolonne of J51044 : Label is "0";
   attribute kolonne of J51043 : Label is "0";
   attribute kolonne of J51042 : Label is "0";
   attribute kolonne of J51041 : Label is "0";
   attribute kolonne of J51040 : Label is "0";
   attribute kolonne of J51039 : Label is "0";
   attribute kolonne of J51038 : Label is "0";
   attribute kolonne of J51037 : Label is "0";
   attribute kolonne of J51036 : Label is "0";
   attribute kolonne of J51035 : Label is "0";
   attribute kolonne of J51034 : Label is "0";
   attribute kolonne of J51033 : Label is "0";
   attribute kolonne of J51032 : Label is "0";
   attribute kolonne of J51031 : Label is "0";
   attribute kolonne of J51030 : Label is "0";
   attribute kolonne of J51029 : Label is "0";
   attribute kolonne of D51003 : Label is "0";
   attribute kolonne of D51002 : Label is "0";
   attribute kolonne of D51001 : Label is "0";

   attribute lager_type : string;
   attribute lager_type of R51046 : Label is "Fremlager";
   attribute lager_type of R51045 : Label is "Fremlager";
   attribute lager_type of R51044 : Label is "Fremlager";
   attribute lager_type of R51043 : Label is "Fremlager";
   attribute lager_type of R51042 : Label is "Fremlager";
   attribute lager_type of R51041 : Label is "Fremlager";
   attribute lager_type of Q51015 : Label is "Fremlager";
   attribute lager_type of Q51014 : Label is "Fremlager";
   attribute lager_type of Q51013 : Label is "Fremlager";
   attribute lager_type of J51049 : Label is "Fremlager";
   attribute lager_type of J51048 : Label is "Fremlager";
   attribute lager_type of J51047 : Label is "Fremlager";
   attribute lager_type of J51046 : Label is "Fremlager";
   attribute lager_type of J51045 : Label is "Fremlager";
   attribute lager_type of J51044 : Label is "Fremlager";
   attribute lager_type of J51043 : Label is "Fremlager";
   attribute lager_type of J51042 : Label is "Fremlager";
   attribute lager_type of J51041 : Label is "Fremlager";
   attribute lager_type of J51040 : Label is "Fremlager";
   attribute lager_type of J51039 : Label is "Fremlager";
   attribute lager_type of J51038 : Label is "Fremlager";
   attribute lager_type of J51037 : Label is "Fremlager";
   attribute lager_type of J51036 : Label is "Fremlager";
   attribute lager_type of J51035 : Label is "Fremlager";
   attribute lager_type of J51034 : Label is "Fremlager";
   attribute lager_type of J51033 : Label is "Fremlager";
   attribute lager_type of J51032 : Label is "Fremlager";
   attribute lager_type of J51031 : Label is "Fremlager";
   attribute lager_type of J51030 : Label is "Fremlager";
   attribute lager_type of J51029 : Label is "Fremlager";
   attribute lager_type of D51003 : Label is "Fremlager";
   attribute lager_type of D51002 : Label is "Fremlager";
   attribute lager_type of D51001 : Label is "Fremlager";

   attribute leverandor : string;
   attribute leverandor of R51043 : Label is "Farnell";
   attribute leverandor of R51042 : Label is "Farnell";
   attribute leverandor of R51041 : Label is "Farnell";
   attribute leverandor of Q51018 : Label is "Farnell";
   attribute leverandor of Q51017 : Label is "Farnell";
   attribute leverandor of Q51016 : Label is "Farnell";
   attribute leverandor of Q51015 : Label is "Farnell";
   attribute leverandor of Q51014 : Label is "Farnell";
   attribute leverandor of Q51013 : Label is "Farnell";
   attribute leverandor of J51028 : Label is "Farnell";
   attribute leverandor of J51008 : Label is "Farnell";
   attribute leverandor of J51007 : Label is "Farnell";
   attribute leverandor of D51003 : Label is "Farnell";
   attribute leverandor of D51002 : Label is "Farnell";
   attribute leverandor of D51001 : Label is "Farnell";

   attribute leverandor_varenr : string;
   attribute leverandor_varenr of R51043 : Label is "2447230";
   attribute leverandor_varenr of R51042 : Label is "2447230";
   attribute leverandor_varenr of R51041 : Label is "2447230";
   attribute leverandor_varenr of Q51018 : Label is "1758073";
   attribute leverandor_varenr of Q51017 : Label is "1758073";
   attribute leverandor_varenr of Q51016 : Label is "1758073";
   attribute leverandor_varenr of Q51015 : Label is "1829184";
   attribute leverandor_varenr of Q51014 : Label is "1829184";
   attribute leverandor_varenr of Q51013 : Label is "1829184";
   attribute leverandor_varenr of J51028 : Label is "1144435";
   attribute leverandor_varenr of J51008 : Label is "1144435";
   attribute leverandor_varenr of J51007 : Label is "1144435";
   attribute leverandor_varenr of D51003 : Label is "8554641";
   attribute leverandor_varenr of D51002 : Label is "8554641";
   attribute leverandor_varenr of D51001 : Label is "8554641";

   attribute navn : string;
   attribute navn of R51046 : Label is "330R";
   attribute navn of R51045 : Label is "330R";
   attribute navn of R51044 : Label is "330R";
   attribute navn of R51043 : Label is "10k";
   attribute navn of R51042 : Label is "10k";
   attribute navn of R51041 : Label is "10k";
   attribute navn of Q51018 : Label is "BSH201";
   attribute navn of Q51017 : Label is "BSH201";
   attribute navn of Q51016 : Label is "BSH201";
   attribute navn of Q51015 : Label is "2N7002";
   attribute navn of Q51014 : Label is "2N7002";
   attribute navn of Q51013 : Label is "2N7002";
   attribute navn of J51049 : Label is "JST 2pin";
   attribute navn of J51048 : Label is "JST 2pin";
   attribute navn of J51047 : Label is "JST 2pin";
   attribute navn of J51046 : Label is "JST 2pin";
   attribute navn of J51045 : Label is "JST 2pin";
   attribute navn of J51044 : Label is "JST 2pin";
   attribute navn of J51043 : Label is "JST 2pin";
   attribute navn of J51042 : Label is "JST 2pin";
   attribute navn of J51041 : Label is "JST 2pin";
   attribute navn of J51040 : Label is "JST 2pin";
   attribute navn of J51039 : Label is "JST 2pin";
   attribute navn of J51038 : Label is "JST 2pin";
   attribute navn of J51037 : Label is "JST 2pin";
   attribute navn of J51036 : Label is "JST 2pin";
   attribute navn of J51035 : Label is "JST 2pin";
   attribute navn of J51034 : Label is "JST 2pin";
   attribute navn of J51033 : Label is "JST 2pin";
   attribute navn of J51032 : Label is "JST 2pin";
   attribute navn of J51031 : Label is "JST 2pin";
   attribute navn of J51030 : Label is "JST 2pin";
   attribute navn of J51029 : Label is "JST 2pin";
   attribute navn of J51028 : Label is "PCI_Express-36P";
   attribute navn of J51008 : Label is "PCI_Express-36P";
   attribute navn of J51007 : Label is "PCI_Express-36P";
   attribute navn of D51003 : Label is "SMD LED Red";
   attribute navn of D51002 : Label is "SMD LED Red";
   attribute navn of D51001 : Label is "SMD LED Red";

   attribute nokkelord : string;
   attribute nokkelord of R51046 : Label is "Resistor Motstand";
   attribute nokkelord of R51045 : Label is "Resistor Motstand";
   attribute nokkelord of R51044 : Label is "Resistor Motstand";
   attribute nokkelord of R51043 : Label is "Resistor Motstand";
   attribute nokkelord of R51042 : Label is "Resistor Motstand";
   attribute nokkelord of R51041 : Label is "Resistor Motstand";
   attribute nokkelord of J51049 : Label is "Connector, Kontakt";
   attribute nokkelord of J51048 : Label is "Connector, Kontakt";
   attribute nokkelord of J51047 : Label is "Connector, Kontakt";
   attribute nokkelord of J51046 : Label is "Connector, Kontakt";
   attribute nokkelord of J51045 : Label is "Connector, Kontakt";
   attribute nokkelord of J51044 : Label is "Connector, Kontakt";
   attribute nokkelord of J51043 : Label is "Connector, Kontakt";
   attribute nokkelord of J51042 : Label is "Connector, Kontakt";
   attribute nokkelord of J51041 : Label is "Connector, Kontakt";
   attribute nokkelord of J51040 : Label is "Connector, Kontakt";
   attribute nokkelord of J51039 : Label is "Connector, Kontakt";
   attribute nokkelord of J51038 : Label is "Connector, Kontakt";
   attribute nokkelord of J51037 : Label is "Connector, Kontakt";
   attribute nokkelord of J51036 : Label is "Connector, Kontakt";
   attribute nokkelord of J51035 : Label is "Connector, Kontakt";
   attribute nokkelord of J51034 : Label is "Connector, Kontakt";
   attribute nokkelord of J51033 : Label is "Connector, Kontakt";
   attribute nokkelord of J51032 : Label is "Connector, Kontakt";
   attribute nokkelord of J51031 : Label is "Connector, Kontakt";
   attribute nokkelord of J51030 : Label is "Connector, Kontakt";
   attribute nokkelord of J51029 : Label is "Connector, Kontakt";
   attribute nokkelord of J51028 : Label is "Card-edge";
   attribute nokkelord of J51008 : Label is "Card-edge";
   attribute nokkelord of J51007 : Label is "Card-edge";
   attribute nokkelord of D51003 : Label is "SMD";
   attribute nokkelord of D51002 : Label is "SMD";
   attribute nokkelord of D51001 : Label is "SMD";

   attribute pakke_opprettet : string;
   attribute pakke_opprettet of R51046 : Label is "08.07.2014 21.15.30";
   attribute pakke_opprettet of R51045 : Label is "08.07.2014 21.15.30";
   attribute pakke_opprettet of R51044 : Label is "08.07.2014 21.15.30";
   attribute pakke_opprettet of R51043 : Label is "08.07.2014 21.15.30";
   attribute pakke_opprettet of R51042 : Label is "08.07.2014 21.15.30";
   attribute pakke_opprettet of R51041 : Label is "08.07.2014 21.15.30";
   attribute pakke_opprettet of Q51018 : Label is "08.07.2014 20.37.25";
   attribute pakke_opprettet of Q51017 : Label is "08.07.2014 20.37.25";
   attribute pakke_opprettet of Q51016 : Label is "08.07.2014 20.37.25";
   attribute pakke_opprettet of Q51015 : Label is "08.07.2014 20.37.25";
   attribute pakke_opprettet of Q51014 : Label is "08.07.2014 20.37.25";
   attribute pakke_opprettet of Q51013 : Label is "08.07.2014 20.37.25";
   attribute pakke_opprettet of J51049 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51048 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51047 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51046 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51045 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51044 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51043 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51042 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51041 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51040 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51039 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51038 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51037 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51036 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51035 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51034 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51033 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51032 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51031 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51030 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51029 : Label is "28.06.2014 18.25.03";
   attribute pakke_opprettet of J51028 : Label is "06.07.2014 17.26.47";
   attribute pakke_opprettet of J51008 : Label is "06.07.2014 17.26.47";
   attribute pakke_opprettet of J51007 : Label is "06.07.2014 17.26.47";
   attribute pakke_opprettet of D51003 : Label is "06.07.2014 18.55.44";
   attribute pakke_opprettet of D51002 : Label is "06.07.2014 18.55.44";
   attribute pakke_opprettet of D51001 : Label is "06.07.2014 18.55.44";

   attribute pakke_opprettet_av : string;
   attribute pakke_opprettet_av of R51046 : Label is "815";
   attribute pakke_opprettet_av of R51045 : Label is "815";
   attribute pakke_opprettet_av of R51044 : Label is "815";
   attribute pakke_opprettet_av of R51043 : Label is "815";
   attribute pakke_opprettet_av of R51042 : Label is "815";
   attribute pakke_opprettet_av of R51041 : Label is "815";
   attribute pakke_opprettet_av of Q51018 : Label is "815";
   attribute pakke_opprettet_av of Q51017 : Label is "815";
   attribute pakke_opprettet_av of Q51016 : Label is "815";
   attribute pakke_opprettet_av of Q51015 : Label is "815";
   attribute pakke_opprettet_av of Q51014 : Label is "815";
   attribute pakke_opprettet_av of Q51013 : Label is "815";
   attribute pakke_opprettet_av of J51049 : Label is "815";
   attribute pakke_opprettet_av of J51048 : Label is "815";
   attribute pakke_opprettet_av of J51047 : Label is "815";
   attribute pakke_opprettet_av of J51046 : Label is "815";
   attribute pakke_opprettet_av of J51045 : Label is "815";
   attribute pakke_opprettet_av of J51044 : Label is "815";
   attribute pakke_opprettet_av of J51043 : Label is "815";
   attribute pakke_opprettet_av of J51042 : Label is "815";
   attribute pakke_opprettet_av of J51041 : Label is "815";
   attribute pakke_opprettet_av of J51040 : Label is "815";
   attribute pakke_opprettet_av of J51039 : Label is "815";
   attribute pakke_opprettet_av of J51038 : Label is "815";
   attribute pakke_opprettet_av of J51037 : Label is "815";
   attribute pakke_opprettet_av of J51036 : Label is "815";
   attribute pakke_opprettet_av of J51035 : Label is "815";
   attribute pakke_opprettet_av of J51034 : Label is "815";
   attribute pakke_opprettet_av of J51033 : Label is "815";
   attribute pakke_opprettet_av of J51032 : Label is "815";
   attribute pakke_opprettet_av of J51031 : Label is "815";
   attribute pakke_opprettet_av of J51030 : Label is "815";
   attribute pakke_opprettet_av of J51029 : Label is "815";
   attribute pakke_opprettet_av of J51028 : Label is "815";
   attribute pakke_opprettet_av of J51008 : Label is "815";
   attribute pakke_opprettet_av of J51007 : Label is "815";
   attribute pakke_opprettet_av of D51003 : Label is "815";
   attribute pakke_opprettet_av of D51002 : Label is "815";
   attribute pakke_opprettet_av of D51001 : Label is "815";

   attribute pakketype : string;
   attribute pakketype of R51046 : Label is "0603";
   attribute pakketype of R51045 : Label is "0603";
   attribute pakketype of R51044 : Label is "0603";
   attribute pakketype of R51043 : Label is "0603";
   attribute pakketype of R51042 : Label is "0603";
   attribute pakketype of R51041 : Label is "0603";
   attribute pakketype of Q51018 : Label is "SOT";
   attribute pakketype of Q51017 : Label is "SOT";
   attribute pakketype of Q51016 : Label is "SOT";
   attribute pakketype of Q51015 : Label is "SMD";
   attribute pakketype of Q51014 : Label is "SMD";
   attribute pakketype of Q51013 : Label is "SMD";
   attribute pakketype of J51049 : Label is "TH";
   attribute pakketype of J51048 : Label is "TH";
   attribute pakketype of J51047 : Label is "TH";
   attribute pakketype of J51046 : Label is "TH";
   attribute pakketype of J51045 : Label is "TH";
   attribute pakketype of J51044 : Label is "TH";
   attribute pakketype of J51043 : Label is "TH";
   attribute pakketype of J51042 : Label is "TH";
   attribute pakketype of J51041 : Label is "TH";
   attribute pakketype of J51040 : Label is "TH";
   attribute pakketype of J51039 : Label is "TH";
   attribute pakketype of J51038 : Label is "TH";
   attribute pakketype of J51037 : Label is "TH";
   attribute pakketype of J51036 : Label is "TH";
   attribute pakketype of J51035 : Label is "TH";
   attribute pakketype of J51034 : Label is "TH";
   attribute pakketype of J51033 : Label is "TH";
   attribute pakketype of J51032 : Label is "TH";
   attribute pakketype of J51031 : Label is "TH";
   attribute pakketype of J51030 : Label is "TH";
   attribute pakketype of J51029 : Label is "TH";
   attribute pakketype of J51028 : Label is "TH";
   attribute pakketype of J51008 : Label is "TH";
   attribute pakketype of J51007 : Label is "TH";
   attribute pakketype of D51003 : Label is "0603";
   attribute pakketype of D51002 : Label is "0603";
   attribute pakketype of D51001 : Label is "0603";

   attribute pris : string;
   attribute pris of R51046 : Label is "0";
   attribute pris of R51045 : Label is "0";
   attribute pris of R51044 : Label is "0";
   attribute pris of R51043 : Label is "0";
   attribute pris of R51042 : Label is "0";
   attribute pris of R51041 : Label is "0";
   attribute pris of Q51018 : Label is "3";
   attribute pris of Q51017 : Label is "3";
   attribute pris of Q51016 : Label is "3";
   attribute pris of Q51015 : Label is "2";
   attribute pris of Q51014 : Label is "2";
   attribute pris of Q51013 : Label is "2";
   attribute pris of J51049 : Label is "2";
   attribute pris of J51048 : Label is "2";
   attribute pris of J51047 : Label is "2";
   attribute pris of J51046 : Label is "2";
   attribute pris of J51045 : Label is "2";
   attribute pris of J51044 : Label is "2";
   attribute pris of J51043 : Label is "2";
   attribute pris of J51042 : Label is "2";
   attribute pris of J51041 : Label is "2";
   attribute pris of J51040 : Label is "2";
   attribute pris of J51039 : Label is "2";
   attribute pris of J51038 : Label is "2";
   attribute pris of J51037 : Label is "2";
   attribute pris of J51036 : Label is "2";
   attribute pris of J51035 : Label is "2";
   attribute pris of J51034 : Label is "2";
   attribute pris of J51033 : Label is "2";
   attribute pris of J51032 : Label is "2";
   attribute pris of J51031 : Label is "2";
   attribute pris of J51030 : Label is "2";
   attribute pris of J51029 : Label is "2";
   attribute pris of J51028 : Label is "16";
   attribute pris of J51008 : Label is "16";
   attribute pris of J51007 : Label is "16";
   attribute pris of D51003 : Label is "1";
   attribute pris of D51002 : Label is "1";
   attribute pris of D51001 : Label is "1";

   attribute produsent : string;
   attribute produsent of R51043 : Label is "Multikomp";
   attribute produsent of R51042 : Label is "Multikomp";
   attribute produsent of R51041 : Label is "Multikomp";
   attribute produsent of Q51018 : Label is "NXP Semiconductors";
   attribute produsent of Q51017 : Label is "NXP Semiconductors";
   attribute produsent of Q51016 : Label is "NXP Semiconductors";
   attribute produsent of J51028 : Label is "FCI";
   attribute produsent of J51008 : Label is "FCI";
   attribute produsent of J51007 : Label is "FCI";
   attribute produsent of D51003 : Label is "Avago";
   attribute produsent of D51002 : Label is "Avago";
   attribute produsent of D51001 : Label is "Avago";

   attribute rad : string;
   attribute rad of R51046 : Label is "-1";
   attribute rad of R51045 : Label is "-1";
   attribute rad of R51044 : Label is "-1";
   attribute rad of R51043 : Label is "-1";
   attribute rad of R51042 : Label is "-1";
   attribute rad of R51041 : Label is "-1";
   attribute rad of Q51015 : Label is "2";
   attribute rad of Q51014 : Label is "2";
   attribute rad of Q51013 : Label is "2";
   attribute rad of J51049 : Label is "3";
   attribute rad of J51048 : Label is "3";
   attribute rad of J51047 : Label is "3";
   attribute rad of J51046 : Label is "3";
   attribute rad of J51045 : Label is "3";
   attribute rad of J51044 : Label is "3";
   attribute rad of J51043 : Label is "3";
   attribute rad of J51042 : Label is "3";
   attribute rad of J51041 : Label is "3";
   attribute rad of J51040 : Label is "3";
   attribute rad of J51039 : Label is "3";
   attribute rad of J51038 : Label is "3";
   attribute rad of J51037 : Label is "3";
   attribute rad of J51036 : Label is "3";
   attribute rad of J51035 : Label is "3";
   attribute rad of J51034 : Label is "3";
   attribute rad of J51033 : Label is "3";
   attribute rad of J51032 : Label is "3";
   attribute rad of J51031 : Label is "3";
   attribute rad of J51030 : Label is "3";
   attribute rad of J51029 : Label is "3";
   attribute rad of D51003 : Label is "0";
   attribute rad of D51002 : Label is "0";
   attribute rad of D51001 : Label is "0";

   attribute rom : string;
   attribute rom of R51046 : Label is "OV";
   attribute rom of R51045 : Label is "OV";
   attribute rom of R51044 : Label is "OV";
   attribute rom of R51043 : Label is "OV";
   attribute rom of R51042 : Label is "OV";
   attribute rom of R51041 : Label is "OV";
   attribute rom of Q51015 : Label is "OV";
   attribute rom of Q51014 : Label is "OV";
   attribute rom of Q51013 : Label is "OV";
   attribute rom of J51049 : Label is "OV";
   attribute rom of J51048 : Label is "OV";
   attribute rom of J51047 : Label is "OV";
   attribute rom of J51046 : Label is "OV";
   attribute rom of J51045 : Label is "OV";
   attribute rom of J51044 : Label is "OV";
   attribute rom of J51043 : Label is "OV";
   attribute rom of J51042 : Label is "OV";
   attribute rom of J51041 : Label is "OV";
   attribute rom of J51040 : Label is "OV";
   attribute rom of J51039 : Label is "OV";
   attribute rom of J51038 : Label is "OV";
   attribute rom of J51037 : Label is "OV";
   attribute rom of J51036 : Label is "OV";
   attribute rom of J51035 : Label is "OV";
   attribute rom of J51034 : Label is "OV";
   attribute rom of J51033 : Label is "OV";
   attribute rom of J51032 : Label is "OV";
   attribute rom of J51031 : Label is "OV";
   attribute rom of J51030 : Label is "OV";
   attribute rom of J51029 : Label is "OV";
   attribute rom of D51003 : Label is "OV";
   attribute rom of D51002 : Label is "OV";
   attribute rom of D51001 : Label is "OV";

   attribute Status : string;
   attribute Status of Q51018 : Label is "New";
   attribute Status of Q51017 : Label is "New";
   attribute Status of Q51016 : Label is "New";

   attribute symbol_opprettet : string;
   attribute symbol_opprettet of R51046 : Label is "08.07.2014 21.16.33";
   attribute symbol_opprettet of R51045 : Label is "08.07.2014 21.16.33";
   attribute symbol_opprettet of R51044 : Label is "08.07.2014 21.16.33";
   attribute symbol_opprettet of R51043 : Label is "08.07.2014 21.16.33";
   attribute symbol_opprettet of R51042 : Label is "08.07.2014 21.16.33";
   attribute symbol_opprettet of R51041 : Label is "08.07.2014 21.16.33";
   attribute symbol_opprettet of Q51018 : Label is "14.09.2016 17.47.57";
   attribute symbol_opprettet of Q51017 : Label is "14.09.2016 17.47.57";
   attribute symbol_opprettet of Q51016 : Label is "14.09.2016 17.47.57";
   attribute symbol_opprettet of Q51015 : Label is "11.07.2014 23.17.04";
   attribute symbol_opprettet of Q51014 : Label is "11.07.2014 23.17.04";
   attribute symbol_opprettet of Q51013 : Label is "11.07.2014 23.17.04";
   attribute symbol_opprettet of J51049 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51048 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51047 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51046 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51045 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51044 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51043 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51042 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51041 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51040 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51039 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51038 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51037 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51036 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51035 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51034 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51033 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51032 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51031 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51030 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51029 : Label is "28.06.2014 15.33.17";
   attribute symbol_opprettet of J51028 : Label is "06.07.2014 17.26.37";
   attribute symbol_opprettet of J51008 : Label is "06.07.2014 17.26.37";
   attribute symbol_opprettet of J51007 : Label is "06.07.2014 17.26.37";
   attribute symbol_opprettet of D51003 : Label is "06.07.2014 18.59.47";
   attribute symbol_opprettet of D51002 : Label is "06.07.2014 18.59.47";
   attribute symbol_opprettet of D51001 : Label is "06.07.2014 18.59.47";

   attribute symbol_opprettet_av : string;
   attribute symbol_opprettet_av of R51046 : Label is "815";
   attribute symbol_opprettet_av of R51045 : Label is "815";
   attribute symbol_opprettet_av of R51044 : Label is "815";
   attribute symbol_opprettet_av of R51043 : Label is "815";
   attribute symbol_opprettet_av of R51042 : Label is "815";
   attribute symbol_opprettet_av of R51041 : Label is "815";
   attribute symbol_opprettet_av of Q51018 : Label is "1150";
   attribute symbol_opprettet_av of Q51017 : Label is "1150";
   attribute symbol_opprettet_av of Q51016 : Label is "1150";
   attribute symbol_opprettet_av of Q51015 : Label is "774";
   attribute symbol_opprettet_av of Q51014 : Label is "774";
   attribute symbol_opprettet_av of Q51013 : Label is "774";
   attribute symbol_opprettet_av of J51049 : Label is "815";
   attribute symbol_opprettet_av of J51048 : Label is "815";
   attribute symbol_opprettet_av of J51047 : Label is "815";
   attribute symbol_opprettet_av of J51046 : Label is "815";
   attribute symbol_opprettet_av of J51045 : Label is "815";
   attribute symbol_opprettet_av of J51044 : Label is "815";
   attribute symbol_opprettet_av of J51043 : Label is "815";
   attribute symbol_opprettet_av of J51042 : Label is "815";
   attribute symbol_opprettet_av of J51041 : Label is "815";
   attribute symbol_opprettet_av of J51040 : Label is "815";
   attribute symbol_opprettet_av of J51039 : Label is "815";
   attribute symbol_opprettet_av of J51038 : Label is "815";
   attribute symbol_opprettet_av of J51037 : Label is "815";
   attribute symbol_opprettet_av of J51036 : Label is "815";
   attribute symbol_opprettet_av of J51035 : Label is "815";
   attribute symbol_opprettet_av of J51034 : Label is "815";
   attribute symbol_opprettet_av of J51033 : Label is "815";
   attribute symbol_opprettet_av of J51032 : Label is "815";
   attribute symbol_opprettet_av of J51031 : Label is "815";
   attribute symbol_opprettet_av of J51030 : Label is "815";
   attribute symbol_opprettet_av of J51029 : Label is "815";
   attribute symbol_opprettet_av of J51028 : Label is "815";
   attribute symbol_opprettet_av of J51008 : Label is "815";
   attribute symbol_opprettet_av of J51007 : Label is "815";
   attribute symbol_opprettet_av of D51003 : Label is "815";
   attribute symbol_opprettet_av of D51002 : Label is "815";
   attribute symbol_opprettet_av of D51001 : Label is "815";

   attribute Verified_by : string;
   attribute Verified_by of Q51018 : Label is "";
   attribute Verified_by of Q51017 : Label is "";
   attribute Verified_by of Q51016 : Label is "";

   attribute Verified_date : string;
   attribute Verified_date of Q51018 : Label is "";
   attribute Verified_date of Q51017 : Label is "";
   attribute Verified_date of Q51016 : Label is "";


Begin
    R51046 : X_2448                                          -- ObjectKind=Part|PrimaryId=R51046|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D51003_1,                           -- ObjectKind=Pin|PrimaryId=R51046-1
        X_2 => PinSignal_Q51018_2                            -- ObjectKind=Pin|PrimaryId=R51046-2
      );

    R51045 : X_2448                                          -- ObjectKind=Part|PrimaryId=R51045|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D51002_1,                           -- ObjectKind=Pin|PrimaryId=R51045-1
        X_2 => PinSignal_Q51017_2                            -- ObjectKind=Pin|PrimaryId=R51045-2
      );

    R51044 : X_2448                                          -- ObjectKind=Part|PrimaryId=R51044|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D51001_1,                           -- ObjectKind=Pin|PrimaryId=R51044-1
        X_2 => PinSignal_Q51016_2                            -- ObjectKind=Pin|PrimaryId=R51044-2
      );

    R51043 : X_2444                                          -- ObjectKind=Part|PrimaryId=R51043|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51028_B1,                          -- ObjectKind=Pin|PrimaryId=R51043-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R51043-2
      );

    R51042 : X_2444                                          -- ObjectKind=Part|PrimaryId=R51042|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51008_B1,                          -- ObjectKind=Pin|PrimaryId=R51042-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R51042-2
      );

    R51041 : X_2444                                          -- ObjectKind=Part|PrimaryId=R51041|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51007_B1,                          -- ObjectKind=Pin|PrimaryId=R51041-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R51041-2
      );

    Q51018 : X_2212                                          -- ObjectKind=Part|PrimaryId=Q51018|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51028_B1,                          -- ObjectKind=Pin|PrimaryId=Q51018-1
        X_2 => PinSignal_Q51018_2,                           -- ObjectKind=Pin|PrimaryId=Q51018-2
        X_3 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=Q51018-3
      );

    Q51017 : X_2212                                          -- ObjectKind=Part|PrimaryId=Q51017|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51008_B1,                          -- ObjectKind=Pin|PrimaryId=Q51017-1
        X_2 => PinSignal_Q51017_2,                           -- ObjectKind=Pin|PrimaryId=Q51017-2
        X_3 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=Q51017-3
      );

    Q51016 : X_2212                                          -- ObjectKind=Part|PrimaryId=Q51016|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51007_B1,                          -- ObjectKind=Pin|PrimaryId=Q51016-1
        X_2 => PinSignal_Q51016_2,                           -- ObjectKind=Pin|PrimaryId=Q51016-2
        X_3 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=Q51016-3
      );

    Q51015 : X_2213                                          -- ObjectKind=Part|PrimaryId=Q51015|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51028_B1,                          -- ObjectKind=Pin|PrimaryId=Q51015-1
        X_2 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=Q51015-2
        X_3 => PinSignal_J51028_A11                          -- ObjectKind=Pin|PrimaryId=Q51015-3
      );

    Q51014 : X_2213                                          -- ObjectKind=Part|PrimaryId=Q51014|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51008_B1,                          -- ObjectKind=Pin|PrimaryId=Q51014-1
        X_2 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=Q51014-2
        X_3 => PinSignal_J51008_A11                          -- ObjectKind=Pin|PrimaryId=Q51014-3
      );

    Q51013 : X_2213                                          -- ObjectKind=Part|PrimaryId=Q51013|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J51007_B1,                          -- ObjectKind=Pin|PrimaryId=Q51013-1
        X_2 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=Q51013-2
        X_3 => PinSignal_J51007_A11                          -- ObjectKind=Pin|PrimaryId=Q51013-3
      );

    J51049 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51049|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51049-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51049-2
      );

    J51048 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51048|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51048-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51048-2
      );

    J51047 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51047|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51047-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51047-2
      );

    J51046 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51046|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51046-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51046-2
      );

    J51045 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51045|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51045-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51045-2
      );

    J51044 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51044|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51044-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51044-2
      );

    J51043 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51043|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51043-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51043-2
      );

    J51042 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51042|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51042-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51042-2
      );

    J51041 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51041|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51041-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51041-2
      );

    J51040 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51040|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51040-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51040-2
      );

    J51039 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51039|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51039-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51039-2
      );

    J51038 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51038|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51038-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51038-2
      );

    J51037 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51037|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51037-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51037-2
      );

    J51036 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51036|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51036-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51036-2
      );

    J51035 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51035|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51035-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51035-2
      );

    J51034 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51034|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51034-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51034-2
      );

    J51033 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51033|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51033-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51033-2
      );

    J51032 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51032|SecondaryId=1
      Port Map
      (
        X_1 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51032-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51032-2
      );

    J51031 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51031|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_AC_S8_L2,                         -- ObjectKind=Pin|PrimaryId=J51031-1
        X_2 => NamedSignal_AC_S8_L1                          -- ObjectKind=Pin|PrimaryId=J51031-2
      );

    J51030 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51030|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_AC_S7_L2,                         -- ObjectKind=Pin|PrimaryId=J51030-1
        X_2 => NamedSignal_AC_S7_L1                          -- ObjectKind=Pin|PrimaryId=J51030-2
      );

    J51029 : X_2227                                          -- ObjectKind=Part|PrimaryId=J51029|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_AC_S6_L2,                         -- ObjectKind=Pin|PrimaryId=J51029-1
        X_2 => NamedSignal_AC_S6_L1                          -- ObjectKind=Pin|PrimaryId=J51029-2
      );

    J51028 : X_2382                                          -- ObjectKind=Part|PrimaryId=J51028|SecondaryId=1
      Port Map
      (
        A1  => PinSignal_J51028_A1,                          -- ObjectKind=Pin|PrimaryId=J51028-A1
        A2  => PinSignal_J51028_A2,                          -- ObjectKind=Pin|PrimaryId=J51028-A2
        A3  => PinSignal_J51028_A3,                          -- ObjectKind=Pin|PrimaryId=J51028-A3
        A4  => PinSignal_J51028_A4,                          -- ObjectKind=Pin|PrimaryId=J51028-A4
        A5  => PinSignal_J51028_A5,                          -- ObjectKind=Pin|PrimaryId=J51028-A5
        A6  => PinSignal_J51028_A6,                          -- ObjectKind=Pin|PrimaryId=J51028-A6
        A7  => PinSignal_J51028_A7,                          -- ObjectKind=Pin|PrimaryId=J51028-A7
        A8  => PinSignal_J51028_A8,                          -- ObjectKind=Pin|PrimaryId=J51028-A8
        A9  => PinSignal_J51028_A9,                          -- ObjectKind=Pin|PrimaryId=J51028-A9
        A10 => PinSignal_J51028_A10,                         -- ObjectKind=Pin|PrimaryId=J51028-A10
        A11 => PinSignal_J51028_A11,                         -- ObjectKind=Pin|PrimaryId=J51028-A11
        A12 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-A12
        A13 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-A13
        A14 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-A14
        A15 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-A15
        A16 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51028-A16
        A17 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51028-A17
        A18 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-A18
        B1  => PinSignal_J51028_B1,                          -- ObjectKind=Pin|PrimaryId=J51028-B1
        B2  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B2
        B3  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B3
        B4  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B4
        B5  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B5
        B6  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B6
        B7  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B7
        B8  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B8
        B9  => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51028-B9
        B11 => NamedSignal_AC_S8_L1,                         -- ObjectKind=Pin|PrimaryId=J51028-B11
        B12 => NamedSignal_AC_S8_L2,                         -- ObjectKind=Pin|PrimaryId=J51028-B12
        B14 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-B14
        B15 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-B15
        B16 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-B16
        B17 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51028-B17
        B18 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51028-B18
      );

    J51008 : X_2382                                          -- ObjectKind=Part|PrimaryId=J51008|SecondaryId=1
      Port Map
      (
        A1  => PinSignal_J51008_A1,                          -- ObjectKind=Pin|PrimaryId=J51008-A1
        A2  => PinSignal_J51008_A2,                          -- ObjectKind=Pin|PrimaryId=J51008-A2
        A3  => PinSignal_J51008_A3,                          -- ObjectKind=Pin|PrimaryId=J51008-A3
        A4  => PinSignal_J51008_A4,                          -- ObjectKind=Pin|PrimaryId=J51008-A4
        A5  => PinSignal_J51008_A5,                          -- ObjectKind=Pin|PrimaryId=J51008-A5
        A6  => PinSignal_J51008_A6,                          -- ObjectKind=Pin|PrimaryId=J51008-A6
        A7  => PinSignal_J51008_A7,                          -- ObjectKind=Pin|PrimaryId=J51008-A7
        A8  => PinSignal_J51008_A8,                          -- ObjectKind=Pin|PrimaryId=J51008-A8
        A9  => PinSignal_J51008_A9,                          -- ObjectKind=Pin|PrimaryId=J51008-A9
        A10 => PinSignal_J51008_A10,                         -- ObjectKind=Pin|PrimaryId=J51008-A10
        A11 => PinSignal_J51008_A11,                         -- ObjectKind=Pin|PrimaryId=J51008-A11
        A12 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-A12
        A13 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-A13
        A14 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-A14
        A15 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-A15
        A16 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51008-A16
        A17 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-A17
        A18 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51008-A18
        B1  => PinSignal_J51008_B1,                          -- ObjectKind=Pin|PrimaryId=J51008-B1
        B2  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B2
        B3  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B3
        B4  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B4
        B5  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B5
        B6  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B6
        B7  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B7
        B8  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B8
        B9  => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51008-B9
        B11 => NamedSignal_AC_S7_L1,                         -- ObjectKind=Pin|PrimaryId=J51008-B11
        B12 => NamedSignal_AC_S7_L2,                         -- ObjectKind=Pin|PrimaryId=J51008-B12
        B14 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-B14
        B15 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-B15
        B16 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-B16
        B17 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51008-B17
        B18 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51008-B18
      );

    J51007 : X_2382                                          -- ObjectKind=Part|PrimaryId=J51007|SecondaryId=1
      Port Map
      (
        A1  => PinSignal_J51007_A1,                          -- ObjectKind=Pin|PrimaryId=J51007-A1
        A2  => PinSignal_J51007_A2,                          -- ObjectKind=Pin|PrimaryId=J51007-A2
        A3  => PinSignal_J51007_A3,                          -- ObjectKind=Pin|PrimaryId=J51007-A3
        A4  => PinSignal_J51007_A4,                          -- ObjectKind=Pin|PrimaryId=J51007-A4
        A5  => PinSignal_J51007_A5,                          -- ObjectKind=Pin|PrimaryId=J51007-A5
        A6  => PinSignal_J51007_A6,                          -- ObjectKind=Pin|PrimaryId=J51007-A6
        A7  => PinSignal_J51007_A7,                          -- ObjectKind=Pin|PrimaryId=J51007-A7
        A8  => PinSignal_J51007_A8,                          -- ObjectKind=Pin|PrimaryId=J51007-A8
        A9  => PinSignal_J51007_A9,                          -- ObjectKind=Pin|PrimaryId=J51007-A9
        A10 => PinSignal_J51007_A10,                         -- ObjectKind=Pin|PrimaryId=J51007-A10
        A11 => PinSignal_J51007_A11,                         -- ObjectKind=Pin|PrimaryId=J51007-A11
        A12 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-A12
        A13 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-A13
        A14 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-A14
        A15 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-A15
        A16 => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-A16
        A17 => PowerSignal_VCC_P5V0,                         -- ObjectKind=Pin|PrimaryId=J51007-A17
        A18 => PowerSignal_VCC_P18V,                         -- ObjectKind=Pin|PrimaryId=J51007-A18
        B1  => PinSignal_J51007_B1,                          -- ObjectKind=Pin|PrimaryId=J51007-B1
        B2  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B2
        B3  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B3
        B4  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B4
        B5  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B5
        B6  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B6
        B7  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B7
        B8  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B8
        B9  => PowerSignal_VCC_EXTRA,                        -- ObjectKind=Pin|PrimaryId=J51007-B9
        B11 => NamedSignal_AC_S6_L1,                         -- ObjectKind=Pin|PrimaryId=J51007-B11
        B12 => NamedSignal_AC_S6_L2,                         -- ObjectKind=Pin|PrimaryId=J51007-B12
        B14 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-B14
        B15 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-B15
        B16 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-B16
        B17 => PowerSignal_GND,                              -- ObjectKind=Pin|PrimaryId=J51007-B17
        B18 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J51007-B18
      );

    D51003 : X_2209                                          -- ObjectKind=Part|PrimaryId=D51003|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D51003_1,                           -- ObjectKind=Pin|PrimaryId=D51003-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D51003-2
      );

    D51002 : X_2209                                          -- ObjectKind=Part|PrimaryId=D51002|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D51002_1,                           -- ObjectKind=Pin|PrimaryId=D51002-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D51002-2
      );

    D51001 : X_2209                                          -- ObjectKind=Part|PrimaryId=D51001|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D51001_1,                           -- ObjectKind=Pin|PrimaryId=D51001-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D51001-2
      );

    -- Signal Assignments
    ---------------------
    BUS_B10              <= PinSignal_J51007_A2; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    BUS_B10              <= PinSignal_J51008_A2; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    BUS_B10              <= PinSignal_J51028_A2; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    BUS_B11              <= PinSignal_J51007_A1; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    BUS_B11              <= PinSignal_J51008_A1; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    BUS_B11              <= PinSignal_J51028_A1; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    BUS_B5               <= PinSignal_J51007_A7; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    BUS_B5               <= PinSignal_J51008_A7; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    BUS_B5               <= PinSignal_J51028_A7; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    BUS_B6               <= PinSignal_J51007_A6; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    BUS_B6               <= PinSignal_J51008_A6; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    BUS_B6               <= PinSignal_J51028_A6; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    BUS_B7               <= PinSignal_J51007_A5; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    BUS_B7               <= PinSignal_J51008_A5; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    BUS_B7               <= PinSignal_J51028_A5; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    BUS_B8               <= PinSignal_J51007_A4; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    BUS_B8               <= PinSignal_J51008_A4; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    BUS_B8               <= PinSignal_J51028_A4; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    BUS_B9               <= PinSignal_J51007_A3; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    BUS_B9               <= PinSignal_J51008_A3; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    BUS_B9               <= PinSignal_J51028_A3; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    BUS_INTERRUPT        <= PinSignal_J51007_A8; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    BUS_INTERRUPT        <= PinSignal_J51008_A8; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    BUS_INTERRUPT        <= PinSignal_J51028_A8; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    BUS_KORT_INNSATT     <= PinSignal_J51007_A11; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    BUS_KORT_INNSATT     <= PinSignal_J51008_A11; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    BUS_KORT_INNSATT     <= PinSignal_J51028_A11; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    BUS_LIMIT            <= PinSignal_J51007_A9; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    BUS_LIMIT            <= PinSignal_J51008_A9; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    BUS_LIMIT            <= PinSignal_J51028_A9; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    BUS_TRIGGER          <= PinSignal_J51007_A10; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    BUS_TRIGGER          <= PinSignal_J51008_A10; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    BUS_TRIGGER          <= PinSignal_J51028_A10; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    PinSignal_J51007_A1  <= BUS_B11; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    PinSignal_J51007_A10 <= BUS_TRIGGER; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    PinSignal_J51007_A11 <= BUS_KORT_INNSATT; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    PinSignal_J51007_A2  <= BUS_B10; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    PinSignal_J51007_A3  <= BUS_B9; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    PinSignal_J51007_A4  <= BUS_B8; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    PinSignal_J51007_A5  <= BUS_B7; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    PinSignal_J51007_A6  <= BUS_B6; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    PinSignal_J51007_A7  <= BUS_B5; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    PinSignal_J51007_A8  <= BUS_INTERRUPT; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    PinSignal_J51007_A9  <= BUS_LIMIT; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    PinSignal_J51008_A1  <= BUS_B11; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    PinSignal_J51008_A10 <= BUS_TRIGGER; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    PinSignal_J51008_A11 <= BUS_KORT_INNSATT; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    PinSignal_J51008_A2  <= BUS_B10; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    PinSignal_J51008_A3  <= BUS_B9; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    PinSignal_J51008_A4  <= BUS_B8; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    PinSignal_J51008_A5  <= BUS_B7; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    PinSignal_J51008_A6  <= BUS_B6; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    PinSignal_J51008_A7  <= BUS_B5; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    PinSignal_J51008_A8  <= BUS_INTERRUPT; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    PinSignal_J51008_A9  <= BUS_LIMIT; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    PinSignal_J51028_A1  <= BUS_B11; -- ObjectKind=Net|PrimaryId=NetJ51028_A1
    PinSignal_J51028_A10 <= BUS_TRIGGER; -- ObjectKind=Net|PrimaryId=NetJ51028_A10
    PinSignal_J51028_A11 <= BUS_KORT_INNSATT; -- ObjectKind=Net|PrimaryId=NetJ51028_A11
    PinSignal_J51028_A2  <= BUS_B10; -- ObjectKind=Net|PrimaryId=NetJ51028_A2
    PinSignal_J51028_A3  <= BUS_B9; -- ObjectKind=Net|PrimaryId=NetJ51028_A3
    PinSignal_J51028_A4  <= BUS_B8; -- ObjectKind=Net|PrimaryId=NetJ51028_A4
    PinSignal_J51028_A5  <= BUS_B7; -- ObjectKind=Net|PrimaryId=NetJ51028_A5
    PinSignal_J51028_A6  <= BUS_B6; -- ObjectKind=Net|PrimaryId=NetJ51028_A6
    PinSignal_J51028_A7  <= BUS_B5; -- ObjectKind=Net|PrimaryId=NetJ51028_A7
    PinSignal_J51028_A8  <= BUS_INTERRUPT; -- ObjectKind=Net|PrimaryId=NetJ51028_A8
    PinSignal_J51028_A9  <= BUS_LIMIT; -- ObjectKind=Net|PrimaryId=NetJ51028_A9
    PowerSignal_GND      <= '0'; -- ObjectKind=Net|PrimaryId=GND

End Structure;
------------------------------------------------------------

