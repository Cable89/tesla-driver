------------------------------------------------------------
-- VHDL TK519_Spenningsvakt
-- 2015 7 5 14 55 24
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 15.0.7.36915
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK519_Spenningsvakt
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK519_Spenningsvakt Is
  attribute MacroCell : boolean;

End TK519_Spenningsvakt;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK519_Spenningsvakt Is


Begin
End Structure;
------------------------------------------------------------

