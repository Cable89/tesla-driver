------------------------------------------------------------
-- VHDL TK520_GDTMINUSTrafo
-- 2015 7 5 14 55 25
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 15.0.7.36915
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK520_GDTMINUSTrafo
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK520_GDTMINUSTrafo Is
  port
  (
    GDT1_1  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT1_1
    GDT1_2  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT1_2
    GDT1_IN : In    STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT1_IN
    GDT2_1  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT2_1
    GDT2_2  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT2_2
    GDT2_IN : In    STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT2_IN
    GDT3_1  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT3_1
    GDT3_2  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT3_2
    GDT4_1  : Out   STD_LOGIC;                               -- ObjectKind=Port|PrimaryId=GDT4_1
    GDT4_2  : Out   STD_LOGIC                                -- ObjectKind=Port|PrimaryId=GDT4_2
  );
  attribute MacroCell : boolean;

End TK520_GDTMINUSTrafo;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK520_GDTMINUSTrafo Is
   Component JST_2pin                                        -- ObjectKind=Part|PrimaryId=J52001|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J52001-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=J52001-2
      );
   End Component;

   Component JST_4pin                                        -- ObjectKind=Part|PrimaryId=J52000|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J52000-1
        X_2 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J52000-2
        X_3 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J52000-3
        X_4 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=J52000-4
      );
   End Component;

   Component SD250MINUS3                                     -- ObjectKind=Part|PrimaryId=T52000|SecondaryId=1
      port
      (
        X_1  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=T52000-1
        X_5  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=T52000-5
        X_6  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=T52000-6
        X_7  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=T52000-7
        X_9  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=T52000-9
        X_10 : inout STD_LOGIC                               -- ObjectKind=Pin|PrimaryId=T52000-10
      );
   End Component;


    Signal PinSignal_J52000_1 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52000_1
    Signal PinSignal_J52000_2 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52000_2
    Signal PinSignal_J52000_3 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52000_3
    Signal PinSignal_J52000_4 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52000_4
    Signal PinSignal_J52002_1 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52002_1
    Signal PinSignal_J52002_2 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52002_2
    Signal PinSignal_J52002_3 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52002_3
    Signal PinSignal_J52002_4 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetJ52002_4

   attribute beskrivelse : string;
   attribute beskrivelse of T52001 : Label is "Dual Gate Drive Transformer";
   attribute beskrivelse of T52000 : Label is "Dual Gate Drive Transformer";

   attribute Database_Table_Name : string;
   attribute Database_Table_Name of T52001 : Label is "altium";
   attribute Database_Table_Name of T52000 : Label is "altium";
   attribute Database_Table_Name of J52002 : Label is "altium";
   attribute Database_Table_Name of J52001 : Label is "altium";
   attribute Database_Table_Name of J52000 : Label is "altium";

   attribute navn : string;
   attribute navn of T52001 : Label is "SD250-3";
   attribute navn of T52000 : Label is "SD250-3";

   attribute nokkelord : string;
   attribute nokkelord of T52001 : Label is "GDT, Tesla";
   attribute nokkelord of T52000 : Label is "GDT, Tesla";

   attribute pakke_opprettet : string;
   attribute pakke_opprettet of T52001 : Label is "28.06.2014 18:37:26";
   attribute pakke_opprettet of T52000 : Label is "28.06.2014 18:37:26";

   attribute pakke_opprettet_av : string;
   attribute pakke_opprettet_av of T52001 : Label is "815";
   attribute pakke_opprettet_av of T52000 : Label is "815";

   attribute pakketype : string;
   attribute pakketype of T52001 : Label is "92";
   attribute pakketype of T52000 : Label is "92";

   attribute pris : string;
   attribute pris of T52001 : Label is "-1";
   attribute pris of T52000 : Label is "-1";

   attribute produsent : string;
   attribute produsent of T52001 : Label is "Coilcraft";
   attribute produsent of T52000 : Label is "Coilcraft";

   attribute symbol_opprettet : string;
   attribute symbol_opprettet of T52001 : Label is "28.06.2014 15:27:34";
   attribute symbol_opprettet of T52000 : Label is "28.06.2014 15:27:34";

   attribute symbol_opprettet_av : string;
   attribute symbol_opprettet_av of T52001 : Label is "815";
   attribute symbol_opprettet_av of T52000 : Label is "815";


Begin
    T52001 : SD250MINUS3                                     -- ObjectKind=Part|PrimaryId=T52001|SecondaryId=1
      Port Map
      (
        X_1  => GDT2_IN,                                     -- ObjectKind=Pin|PrimaryId=T52001-1
        X_5  => GDT1_IN,                                     -- ObjectKind=Pin|PrimaryId=T52001-5
        X_6  => PinSignal_J52002_1,                          -- ObjectKind=Pin|PrimaryId=T52001-6
        X_7  => PinSignal_J52002_2,                          -- ObjectKind=Pin|PrimaryId=T52001-7
        X_9  => PinSignal_J52002_3,                          -- ObjectKind=Pin|PrimaryId=T52001-9
        X_10 => PinSignal_J52002_4                           -- ObjectKind=Pin|PrimaryId=T52001-10
      );

    T52000 : SD250MINUS3                                     -- ObjectKind=Part|PrimaryId=T52000|SecondaryId=1
      Port Map
      (
        X_1  => GDT1_IN,                                     -- ObjectKind=Pin|PrimaryId=T52000-1
        X_5  => GDT2_IN,                                     -- ObjectKind=Pin|PrimaryId=T52000-5
        X_6  => PinSignal_J52000_1,                          -- ObjectKind=Pin|PrimaryId=T52000-6
        X_7  => PinSignal_J52000_2,                          -- ObjectKind=Pin|PrimaryId=T52000-7
        X_9  => PinSignal_J52000_3,                          -- ObjectKind=Pin|PrimaryId=T52000-9
        X_10 => PinSignal_J52000_4                           -- ObjectKind=Pin|PrimaryId=T52000-10
      );

    J52002 : JST_4pin                                        -- ObjectKind=Part|PrimaryId=J52002|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J52002_1,                           -- ObjectKind=Pin|PrimaryId=J52002-1
        X_2 => PinSignal_J52002_2,                           -- ObjectKind=Pin|PrimaryId=J52002-2
        X_3 => PinSignal_J52002_3,                           -- ObjectKind=Pin|PrimaryId=J52002-3
        X_4 => PinSignal_J52002_4                            -- ObjectKind=Pin|PrimaryId=J52002-4
      );

    J52001 : JST_2pin                                        -- ObjectKind=Part|PrimaryId=J52001|SecondaryId=1
      Port Map
      (
        X_1 => GDT1_IN,                                      -- ObjectKind=Pin|PrimaryId=J52001-1
        X_2 => GDT2_IN                                       -- ObjectKind=Pin|PrimaryId=J52001-2
      );

    J52000 : JST_4pin                                        -- ObjectKind=Part|PrimaryId=J52000|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_J52000_1,                           -- ObjectKind=Pin|PrimaryId=J52000-1
        X_2 => PinSignal_J52000_2,                           -- ObjectKind=Pin|PrimaryId=J52000-2
        X_3 => PinSignal_J52000_3,                           -- ObjectKind=Pin|PrimaryId=J52000-3
        X_4 => PinSignal_J52000_4                            -- ObjectKind=Pin|PrimaryId=J52000-4
      );

    -- Signal Assignments
    ---------------------
    GDT1_1             <= PinSignal_J52000_1; -- ObjectKind=Net|PrimaryId=NetJ52000_1
    GDT1_2             <= PinSignal_J52002_1; -- ObjectKind=Net|PrimaryId=NetJ52002_1
    GDT2_1             <= PinSignal_J52000_2; -- ObjectKind=Net|PrimaryId=NetJ52000_2
    GDT2_2             <= PinSignal_J52002_2; -- ObjectKind=Net|PrimaryId=NetJ52002_2
    GDT3_1             <= PinSignal_J52000_3; -- ObjectKind=Net|PrimaryId=NetJ52000_3
    GDT3_2             <= PinSignal_J52002_3; -- ObjectKind=Net|PrimaryId=NetJ52002_3
    GDT4_1             <= PinSignal_J52000_4; -- ObjectKind=Net|PrimaryId=NetJ52000_4
    GDT4_2             <= PinSignal_J52002_4; -- ObjectKind=Net|PrimaryId=NetJ52002_4
    PinSignal_J52000_1 <= GDT1_1; -- ObjectKind=Net|PrimaryId=NetJ52000_1
    PinSignal_J52000_2 <= GDT2_1; -- ObjectKind=Net|PrimaryId=NetJ52000_2
    PinSignal_J52000_3 <= GDT3_1; -- ObjectKind=Net|PrimaryId=NetJ52000_3
    PinSignal_J52000_4 <= GDT4_1; -- ObjectKind=Net|PrimaryId=NetJ52000_4
    PinSignal_J52002_1 <= GDT1_2; -- ObjectKind=Net|PrimaryId=NetJ52002_1
    PinSignal_J52002_2 <= GDT2_2; -- ObjectKind=Net|PrimaryId=NetJ52002_2
    PinSignal_J52002_3 <= GDT3_2; -- ObjectKind=Net|PrimaryId=NetJ52002_3
    PinSignal_J52002_4 <= GDT4_2; -- ObjectKind=Net|PrimaryId=NetJ52002_4

End Structure;
------------------------------------------------------------

