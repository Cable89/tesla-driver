------------------------------------------------------------
-- VHDL TK530_Kraftbakplan
-- 2014 7 12 23 24 5
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.11.33708
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK530_Kraftbakplan
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK530_Kraftbakplan Is
  port
  (
    GDT1_1    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT1_1
    GDT1_2    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT1_2
    GDT2_1    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT2_1
    GDT2_2    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT2_2
    GDT3_1    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT3_1
    GDT3_2    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT3_2
    GDT4_1    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT4_1
    GDT4_2    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GDT4_2
    GND_HV    : In    STD_LOGIC;                             -- ObjectKind=Port|PrimaryId=GND_HV
    VCC_P18V0 : In    STD_LOGIC                              -- ObjectKind=Port|PrimaryId=VCC_P18V0
  );
  attribute MacroCell : boolean;

End TK530_Kraftbakplan;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK530_Kraftbakplan Is


Begin
End Structure;
------------------------------------------------------------

