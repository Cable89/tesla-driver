------------------------------------------------------------
-- VHDL TK532_Utgangskondensator
-- 2014 7 5 19 58 31
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2004 Altium Limited"
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK532_Utgangskondensator
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK532_Utgangskondensator Is
  attribute MacroCell : boolean;

End TK532_Utgangskondensator;
------------------------------------------------------------

------------------------------------------------------------
architecture structure of TK532_Utgangskondensator is


begin
end structure;
------------------------------------------------------------

