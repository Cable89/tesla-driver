------------------------------------------------------------
-- VHDL TK516_EKSTRAMINUSPSU
-- 2016 1 26 18 15 21
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.0.5.271
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK516_EKSTRAMINUSPSU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK516_EKSTRAMINUSPSU Is
  attribute MacroCell : boolean;

End TK516_EKSTRAMINUSPSU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK516_EKSTRAMINUSPSU Is


Begin
End Structure;
------------------------------------------------------------

