------------------------------------------------------------
-- VHDL TK540_Frontpanel
-- 2016 4 30 0 12 25
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.0.5.271
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK540_Frontpanel
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK540_Frontpanel Is
  attribute MacroCell : boolean;

End TK540_Frontpanel;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK540_Frontpanel Is
   Component TK502_Frontpanel_LEDs                           -- ObjectKind=Sheet Symbol|PrimaryId=LEDs
   End Component;



Begin
    LEDs : TK502_Frontpanel_LEDs                             -- ObjectKind=Sheet Symbol|PrimaryId=LEDs
;

End Structure;
------------------------------------------------------------

