------------------------------------------------------------
-- VHDL TK532_Utgangskondensator
-- 2014 7 12 21 38 42
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK532_Utgangskondensator
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK532_Utgangskondensator Is
  attribute MacroCell : boolean;

End TK532_Utgangskondensator;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK532_Utgangskondensator Is


Begin
End Structure;
------------------------------------------------------------

