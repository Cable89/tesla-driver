------------------------------------------------------------
-- VHDL TK517_P5V0MINUSPSU
-- 2016 9 23 13 35 52
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.0.5.271
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK517_P5V0MINUSPSU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK517_P5V0MINUSPSU Is
  attribute MacroCell : boolean;

End TK517_P5V0MINUSPSU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK517_P5V0MINUSPSU Is


Begin
End Structure;
------------------------------------------------------------

