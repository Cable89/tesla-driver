------------------------------------------------------------
-- VHDL TK517_P5V0MINUSPSU
-- 2016 4 28 20 30 5
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 15.0.15.41991
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK517_P5V0MINUSPSU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK517_P5V0MINUSPSU Is
  attribute MacroCell : boolean;

End TK517_P5V0MINUSPSU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK517_P5V0MINUSPSU Is


Begin
End Structure;
------------------------------------------------------------

