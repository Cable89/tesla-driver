------------------------------------------------------------
-- VHDL TK519_Spenningsvakt
-- 2014 7 6 17 49 12
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.11.33708
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK519_Spenningsvakt
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK519_Spenningsvakt Is
  attribute MacroCell : boolean;

End TK519_Spenningsvakt;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK519_Spenningsvakt Is


Begin
End Structure;
------------------------------------------------------------

