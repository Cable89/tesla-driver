------------------------------------------------------------
-- VHDL TK502_Frontpanel_LEDs
-- 2016 4 28 20 30 6
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 15.0.15.41991
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK502_Frontpanel_LEDs
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK502_Frontpanel_LEDs Is
  attribute MacroCell : boolean;

End TK502_Frontpanel_LEDs;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK502_Frontpanel_LEDs Is
   Component X_2076                                          -- ObjectKind=Part|PrimaryId=D50200|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=D50200-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=D50200-2
      );
   End Component;

   Component X_2226                                          -- ObjectKind=Part|PrimaryId=J50200|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J50200-1
        X_2 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=J50200-2
        X_3 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=J50200-3
      );
   End Component;

   Component X_2384                                          -- ObjectKind=Part|PrimaryId=R50200|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=R50200-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=R50200-2
      );
   End Component;

   Component X_2390                                          -- ObjectKind=Part|PrimaryId=J50206|SecondaryId=1
      port
      (
        X_1  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-1
        X_2  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-2
        X_3  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-3
        X_4  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-4
        X_5  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-5
        X_6  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-6
        X_7  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-7
        X_8  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-8
        X_9  : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-9
        X_10 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-10
        X_11 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-11
        X_12 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-12
        X_13 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-13
        X_14 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-14
        X_15 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-15
        X_16 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-16
        X_17 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-17
        X_18 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-18
        X_19 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-19
        X_20 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-20
        X_21 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-21
        X_22 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-22
        X_23 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-23
        X_24 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-24
        X_25 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-25
        X_26 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-26
        X_27 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-27
        X_28 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-28
        X_29 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-29
        X_30 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-30
        X_31 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-31
        X_32 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-32
        X_33 : inout STD_LOGIC;                              -- ObjectKind=Pin|PrimaryId=J50206-33
        X_34 : inout STD_LOGIC                               -- ObjectKind=Pin|PrimaryId=J50206-34
      );
   End Component;

   Component X_2448                                          -- ObjectKind=Part|PrimaryId=R50202|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=R50202-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=R50202-2
      );
   End Component;

   Component X_3597                                          -- ObjectKind=Part|PrimaryId=D50201|SecondaryId=1
      port
      (
        X_1 : inout STD_LOGIC;                               -- ObjectKind=Pin|PrimaryId=D50201-1
        X_2 : inout STD_LOGIC                                -- ObjectKind=Pin|PrimaryId=D50201-2
      );
   End Component;


    Signal NamedSignal_0_FE     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=0_FE
    Signal NamedSignal_0_INT    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=0_INT
    Signal NamedSignal_0_KI     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=0_KI
    Signal NamedSignal_0_KNP    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=0_KNP
    Signal NamedSignal_0_ST     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=0_ST
    Signal NamedSignal_1_FE     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=1_FE
    Signal NamedSignal_1_INT    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=1_INT
    Signal NamedSignal_1_KI     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=1_KI
    Signal NamedSignal_1_KNP    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=1_KNP
    Signal NamedSignal_1_ST     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=1_ST
    Signal NamedSignal_2_FE     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=2_FE
    Signal NamedSignal_2_INT    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=2_INT
    Signal NamedSignal_2_KI     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=2_KI
    Signal NamedSignal_2_KNP    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=2_KNP
    Signal NamedSignal_2_ST     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=2_ST
    Signal NamedSignal_3_FE     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=3_FE
    Signal NamedSignal_3_INT    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=3_INT
    Signal NamedSignal_3_KI     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=3_KI
    Signal NamedSignal_3_KNP    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=3_KNP
    Signal NamedSignal_3_ST     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=3_ST
    Signal NamedSignal_4_FE     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=4_FE
    Signal NamedSignal_4_INT    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=4_INT
    Signal NamedSignal_4_KI     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=4_KI
    Signal NamedSignal_4_KNP    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=4_KNP
    Signal NamedSignal_4_ST     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=4_ST
    Signal NamedSignal_5_FE     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=5_FE
    Signal NamedSignal_5_INT    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=5_INT
    Signal NamedSignal_5_KI     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=5_KI
    Signal NamedSignal_5_KNP    : STD_LOGIC; -- ObjectKind=Net|PrimaryId=5_KNP
    Signal NamedSignal_5_ST     : STD_LOGIC; -- ObjectKind=Net|PrimaryId=5_ST
    Signal PinSignal_D50200_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50200_1
    Signal PinSignal_D50201_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50201_1
    Signal PinSignal_D50202_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50202_1
    Signal PinSignal_D50203_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50203_1
    Signal PinSignal_D50204_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50204_1
    Signal PinSignal_D50205_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50205_1
    Signal PinSignal_D50206_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50206_1
    Signal PinSignal_D50207_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50207_1
    Signal PinSignal_D50208_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50208_1
    Signal PinSignal_D50209_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50209_1
    Signal PinSignal_D50210_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50210_1
    Signal PinSignal_D50211_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50211_1
    Signal PinSignal_D50212_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50212_1
    Signal PinSignal_D50213_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50213_1
    Signal PinSignal_D50214_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50214_1
    Signal PinSignal_D50215_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50215_1
    Signal PinSignal_D50216_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50216_1
    Signal PinSignal_D50217_1   : STD_LOGIC; -- ObjectKind=Net|PrimaryId=NetD50217_1
    Signal PowerSignal_GND      : STD_LOGIC; -- ObjectKind=Net|PrimaryId=GND
    Signal PowerSignal_VCC_P5V0 : STD_LOGIC; -- ObjectKind=Net|PrimaryId=VCC_P5V0

   attribute antall : string;
   attribute antall of R50223 : Label is "100";
   attribute antall of R50222 : Label is "100";
   attribute antall of R50221 : Label is "100";
   attribute antall of R50220 : Label is "100";
   attribute antall of R50219 : Label is "100";
   attribute antall of R50218 : Label is "100";
   attribute antall of R50217 : Label is "100";
   attribute antall of R50216 : Label is "100";
   attribute antall of R50215 : Label is "100";
   attribute antall of R50214 : Label is "100";
   attribute antall of R50213 : Label is "100";
   attribute antall of R50212 : Label is "100";
   attribute antall of R50211 : Label is "100";
   attribute antall of R50210 : Label is "100";
   attribute antall of R50209 : Label is "100";
   attribute antall of R50208 : Label is "100";
   attribute antall of R50207 : Label is "100";
   attribute antall of R50206 : Label is "100";
   attribute antall of R50205 : Label is "100";
   attribute antall of R50204 : Label is "100";
   attribute antall of R50203 : Label is "100";
   attribute antall of R50202 : Label is "100";
   attribute antall of R50201 : Label is "100";
   attribute antall of R50200 : Label is "100";

   attribute beskrivelse : string;
   attribute beskrivelse of D50217 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50216 : Label is "LED, Red, 5mm, 643 nm, 1.8 V, 20 mA, 400 mcd";
   attribute beskrivelse of D50215 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50214 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50213 : Label is "LED, Red, 5mm, 643 nm, 1.8 V, 20 mA, 400 mcd";
   attribute beskrivelse of D50212 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50211 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50210 : Label is "LED, Red, 5mm, 643 nm, 1.8 V, 20 mA, 400 mcd";
   attribute beskrivelse of D50209 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50208 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50207 : Label is "LED, Red, 5mm, 643 nm, 1.8 V, 20 mA, 400 mcd";
   attribute beskrivelse of D50206 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50205 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50204 : Label is "LED, Red, 5mm, 643 nm, 1.8 V, 20 mA, 400 mcd";
   attribute beskrivelse of D50203 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50202 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";
   attribute beskrivelse of D50201 : Label is "LED, Red, 5mm, 643 nm, 1.8 V, 20 mA, 400 mcd";
   attribute beskrivelse of D50200 : Label is "LED, Green, 5mm, 572 nm, 2.1 V, 20 mA, 150 mcd";

   attribute Database_Table_Name : string;
   attribute Database_Table_Name of R50223 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50222 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50221 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50220 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50219 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50218 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50217 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50216 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50215 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50214 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50213 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50212 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50211 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50210 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50209 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50208 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50207 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50206 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50205 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50204 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50203 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50202 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50201 : Label is "altium_Motstander";
   attribute Database_Table_Name of R50200 : Label is "altium_Motstander";
   attribute Database_Table_Name of J50206 : Label is "altium";
   attribute Database_Table_Name of J50205 : Label is "altium";
   attribute Database_Table_Name of J50204 : Label is "altium";
   attribute Database_Table_Name of J50203 : Label is "altium";
   attribute Database_Table_Name of J50202 : Label is "altium";
   attribute Database_Table_Name of J50201 : Label is "altium";
   attribute Database_Table_Name of J50200 : Label is "altium";
   attribute Database_Table_Name of D50217 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50216 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50215 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50214 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50213 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50212 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50211 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50210 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50209 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50208 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50207 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50206 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50205 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50204 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50203 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50202 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50201 : Label is "altium_Dioder";
   attribute Database_Table_Name of D50200 : Label is "altium_Dioder";

   attribute dybde : string;
   attribute dybde of R50223 : Label is "36";
   attribute dybde of R50222 : Label is "36";
   attribute dybde of R50221 : Label is "36";
   attribute dybde of R50220 : Label is "36";
   attribute dybde of R50219 : Label is "36";
   attribute dybde of R50218 : Label is "36";
   attribute dybde of R50217 : Label is "96";
   attribute dybde of R50216 : Label is "96";
   attribute dybde of R50215 : Label is "36";
   attribute dybde of R50214 : Label is "36";
   attribute dybde of R50213 : Label is "36";
   attribute dybde of R50212 : Label is "36";
   attribute dybde of R50211 : Label is "36";
   attribute dybde of R50210 : Label is "36";
   attribute dybde of R50209 : Label is "96";
   attribute dybde of R50208 : Label is "96";
   attribute dybde of R50207 : Label is "36";
   attribute dybde of R50206 : Label is "36";
   attribute dybde of R50205 : Label is "36";
   attribute dybde of R50204 : Label is "36";
   attribute dybde of R50203 : Label is "36";
   attribute dybde of R50202 : Label is "36";
   attribute dybde of R50201 : Label is "96";
   attribute dybde of R50200 : Label is "96";

   attribute hylle : string;
   attribute hylle of R50223 : Label is "6";
   attribute hylle of R50222 : Label is "6";
   attribute hylle of R50221 : Label is "6";
   attribute hylle of R50220 : Label is "6";
   attribute hylle of R50219 : Label is "6";
   attribute hylle of R50218 : Label is "6";
   attribute hylle of R50217 : Label is "6";
   attribute hylle of R50216 : Label is "6";
   attribute hylle of R50215 : Label is "6";
   attribute hylle of R50214 : Label is "6";
   attribute hylle of R50213 : Label is "6";
   attribute hylle of R50212 : Label is "6";
   attribute hylle of R50211 : Label is "6";
   attribute hylle of R50210 : Label is "6";
   attribute hylle of R50209 : Label is "6";
   attribute hylle of R50208 : Label is "6";
   attribute hylle of R50207 : Label is "6";
   attribute hylle of R50206 : Label is "6";
   attribute hylle of R50205 : Label is "6";
   attribute hylle of R50204 : Label is "6";
   attribute hylle of R50203 : Label is "6";
   attribute hylle of R50202 : Label is "6";
   attribute hylle of R50201 : Label is "6";
   attribute hylle of R50200 : Label is "6";

   attribute id : string;
   attribute id of R50223 : Label is "2448";
   attribute id of R50222 : Label is "2448";
   attribute id of R50221 : Label is "2448";
   attribute id of R50220 : Label is "2448";
   attribute id of R50219 : Label is "2448";
   attribute id of R50218 : Label is "2448";
   attribute id of R50217 : Label is "2384";
   attribute id of R50216 : Label is "2384";
   attribute id of R50215 : Label is "2448";
   attribute id of R50214 : Label is "2448";
   attribute id of R50213 : Label is "2448";
   attribute id of R50212 : Label is "2448";
   attribute id of R50211 : Label is "2448";
   attribute id of R50210 : Label is "2448";
   attribute id of R50209 : Label is "2384";
   attribute id of R50208 : Label is "2384";
   attribute id of R50207 : Label is "2448";
   attribute id of R50206 : Label is "2448";
   attribute id of R50205 : Label is "2448";
   attribute id of R50204 : Label is "2448";
   attribute id of R50203 : Label is "2448";
   attribute id of R50202 : Label is "2448";
   attribute id of R50201 : Label is "2384";
   attribute id of R50200 : Label is "2384";
   attribute id of J50206 : Label is "2390";
   attribute id of J50205 : Label is "2226";
   attribute id of J50204 : Label is "2226";
   attribute id of J50203 : Label is "2226";
   attribute id of J50202 : Label is "2226";
   attribute id of J50201 : Label is "2226";
   attribute id of J50200 : Label is "2226";
   attribute id of D50217 : Label is "2076";
   attribute id of D50216 : Label is "3597";
   attribute id of D50215 : Label is "2076";
   attribute id of D50214 : Label is "2076";
   attribute id of D50213 : Label is "3597";
   attribute id of D50212 : Label is "2076";
   attribute id of D50211 : Label is "2076";
   attribute id of D50210 : Label is "3597";
   attribute id of D50209 : Label is "2076";
   attribute id of D50208 : Label is "2076";
   attribute id of D50207 : Label is "3597";
   attribute id of D50206 : Label is "2076";
   attribute id of D50205 : Label is "2076";
   attribute id of D50204 : Label is "3597";
   attribute id of D50203 : Label is "2076";
   attribute id of D50202 : Label is "2076";
   attribute id of D50201 : Label is "3597";
   attribute id of D50200 : Label is "2076";

   attribute kolonne : string;
   attribute kolonne of R50223 : Label is "0";
   attribute kolonne of R50222 : Label is "0";
   attribute kolonne of R50221 : Label is "0";
   attribute kolonne of R50220 : Label is "0";
   attribute kolonne of R50219 : Label is "0";
   attribute kolonne of R50218 : Label is "0";
   attribute kolonne of R50217 : Label is "0";
   attribute kolonne of R50216 : Label is "0";
   attribute kolonne of R50215 : Label is "0";
   attribute kolonne of R50214 : Label is "0";
   attribute kolonne of R50213 : Label is "0";
   attribute kolonne of R50212 : Label is "0";
   attribute kolonne of R50211 : Label is "0";
   attribute kolonne of R50210 : Label is "0";
   attribute kolonne of R50209 : Label is "0";
   attribute kolonne of R50208 : Label is "0";
   attribute kolonne of R50207 : Label is "0";
   attribute kolonne of R50206 : Label is "0";
   attribute kolonne of R50205 : Label is "0";
   attribute kolonne of R50204 : Label is "0";
   attribute kolonne of R50203 : Label is "0";
   attribute kolonne of R50202 : Label is "0";
   attribute kolonne of R50201 : Label is "0";
   attribute kolonne of R50200 : Label is "0";

   attribute lager_type : string;
   attribute lager_type of R50223 : Label is "Fremlager";
   attribute lager_type of R50222 : Label is "Fremlager";
   attribute lager_type of R50221 : Label is "Fremlager";
   attribute lager_type of R50220 : Label is "Fremlager";
   attribute lager_type of R50219 : Label is "Fremlager";
   attribute lager_type of R50218 : Label is "Fremlager";
   attribute lager_type of R50217 : Label is "Fremlager";
   attribute lager_type of R50216 : Label is "Fremlager";
   attribute lager_type of R50215 : Label is "Fremlager";
   attribute lager_type of R50214 : Label is "Fremlager";
   attribute lager_type of R50213 : Label is "Fremlager";
   attribute lager_type of R50212 : Label is "Fremlager";
   attribute lager_type of R50211 : Label is "Fremlager";
   attribute lager_type of R50210 : Label is "Fremlager";
   attribute lager_type of R50209 : Label is "Fremlager";
   attribute lager_type of R50208 : Label is "Fremlager";
   attribute lager_type of R50207 : Label is "Fremlager";
   attribute lager_type of R50206 : Label is "Fremlager";
   attribute lager_type of R50205 : Label is "Fremlager";
   attribute lager_type of R50204 : Label is "Fremlager";
   attribute lager_type of R50203 : Label is "Fremlager";
   attribute lager_type of R50202 : Label is "Fremlager";
   attribute lager_type of R50201 : Label is "Fremlager";
   attribute lager_type of R50200 : Label is "Fremlager";

   attribute leverandor : string;
   attribute leverandor of D50217 : Label is "Farnell";
   attribute leverandor of D50216 : Label is "Farnell";
   attribute leverandor of D50215 : Label is "Farnell";
   attribute leverandor of D50214 : Label is "Farnell";
   attribute leverandor of D50213 : Label is "Farnell";
   attribute leverandor of D50212 : Label is "Farnell";
   attribute leverandor of D50211 : Label is "Farnell";
   attribute leverandor of D50210 : Label is "Farnell";
   attribute leverandor of D50209 : Label is "Farnell";
   attribute leverandor of D50208 : Label is "Farnell";
   attribute leverandor of D50207 : Label is "Farnell";
   attribute leverandor of D50206 : Label is "Farnell";
   attribute leverandor of D50205 : Label is "Farnell";
   attribute leverandor of D50204 : Label is "Farnell";
   attribute leverandor of D50203 : Label is "Farnell";
   attribute leverandor of D50202 : Label is "Farnell";
   attribute leverandor of D50201 : Label is "Farnell";
   attribute leverandor of D50200 : Label is "Farnell";

   attribute leverandor_varenr : string;
   attribute leverandor_varenr of D50217 : Label is "2112108";
   attribute leverandor_varenr of D50216 : Label is "2112111";
   attribute leverandor_varenr of D50215 : Label is "2112108";
   attribute leverandor_varenr of D50214 : Label is "2112108";
   attribute leverandor_varenr of D50213 : Label is "2112111";
   attribute leverandor_varenr of D50212 : Label is "2112108";
   attribute leverandor_varenr of D50211 : Label is "2112108";
   attribute leverandor_varenr of D50210 : Label is "2112111";
   attribute leverandor_varenr of D50209 : Label is "2112108";
   attribute leverandor_varenr of D50208 : Label is "2112108";
   attribute leverandor_varenr of D50207 : Label is "2112111";
   attribute leverandor_varenr of D50206 : Label is "2112108";
   attribute leverandor_varenr of D50205 : Label is "2112108";
   attribute leverandor_varenr of D50204 : Label is "2112111";
   attribute leverandor_varenr of D50203 : Label is "2112108";
   attribute leverandor_varenr of D50202 : Label is "2112108";
   attribute leverandor_varenr of D50201 : Label is "2112111";
   attribute leverandor_varenr of D50200 : Label is "2112108";

   attribute navn : string;
   attribute navn of R50223 : Label is "330R";
   attribute navn of R50222 : Label is "330R";
   attribute navn of R50221 : Label is "330R";
   attribute navn of R50220 : Label is "330R";
   attribute navn of R50219 : Label is "330R";
   attribute navn of R50218 : Label is "330R";
   attribute navn of R50217 : Label is "100k";
   attribute navn of R50216 : Label is "100k";
   attribute navn of R50215 : Label is "330R";
   attribute navn of R50214 : Label is "330R";
   attribute navn of R50213 : Label is "330R";
   attribute navn of R50212 : Label is "330R";
   attribute navn of R50211 : Label is "330R";
   attribute navn of R50210 : Label is "330R";
   attribute navn of R50209 : Label is "100k";
   attribute navn of R50208 : Label is "100k";
   attribute navn of R50207 : Label is "330R";
   attribute navn of R50206 : Label is "330R";
   attribute navn of R50205 : Label is "330R";
   attribute navn of R50204 : Label is "330R";
   attribute navn of R50203 : Label is "330R";
   attribute navn of R50202 : Label is "330R";
   attribute navn of R50201 : Label is "100k";
   attribute navn of R50200 : Label is "100k";
   attribute navn of J50206 : Label is "Header Shrouded 2X17P";
   attribute navn of J50205 : Label is "JST 3pin";
   attribute navn of J50204 : Label is "JST 3pin";
   attribute navn of J50203 : Label is "JST 3pin";
   attribute navn of J50202 : Label is "JST 3pin";
   attribute navn of J50201 : Label is "JST 3pin";
   attribute navn of J50200 : Label is "JST 3pin";
   attribute navn of D50217 : Label is "Gr�nn LED 5mm";
   attribute navn of D50216 : Label is "R�d LED 5mm";
   attribute navn of D50215 : Label is "Gr�nn LED 5mm";
   attribute navn of D50214 : Label is "Gr�nn LED 5mm";
   attribute navn of D50213 : Label is "R�d LED 5mm";
   attribute navn of D50212 : Label is "Gr�nn LED 5mm";
   attribute navn of D50211 : Label is "Gr�nn LED 5mm";
   attribute navn of D50210 : Label is "R�d LED 5mm";
   attribute navn of D50209 : Label is "Gr�nn LED 5mm";
   attribute navn of D50208 : Label is "Gr�nn LED 5mm";
   attribute navn of D50207 : Label is "R�d LED 5mm";
   attribute navn of D50206 : Label is "Gr�nn LED 5mm";
   attribute navn of D50205 : Label is "Gr�nn LED 5mm";
   attribute navn of D50204 : Label is "R�d LED 5mm";
   attribute navn of D50203 : Label is "Gr�nn LED 5mm";
   attribute navn of D50202 : Label is "Gr�nn LED 5mm";
   attribute navn of D50201 : Label is "R�d LED 5mm";
   attribute navn of D50200 : Label is "Gr�nn LED 5mm";

   attribute nokkelord : string;
   attribute nokkelord of R50223 : Label is "Resistor Motstand";
   attribute nokkelord of R50222 : Label is "Resistor Motstand";
   attribute nokkelord of R50221 : Label is "Resistor Motstand";
   attribute nokkelord of R50220 : Label is "Resistor Motstand";
   attribute nokkelord of R50219 : Label is "Resistor Motstand";
   attribute nokkelord of R50218 : Label is "Resistor Motstand";
   attribute nokkelord of R50217 : Label is "Resistor";
   attribute nokkelord of R50216 : Label is "Resistor";
   attribute nokkelord of R50215 : Label is "Resistor Motstand";
   attribute nokkelord of R50214 : Label is "Resistor Motstand";
   attribute nokkelord of R50213 : Label is "Resistor Motstand";
   attribute nokkelord of R50212 : Label is "Resistor Motstand";
   attribute nokkelord of R50211 : Label is "Resistor Motstand";
   attribute nokkelord of R50210 : Label is "Resistor Motstand";
   attribute nokkelord of R50209 : Label is "Resistor";
   attribute nokkelord of R50208 : Label is "Resistor";
   attribute nokkelord of R50207 : Label is "Resistor Motstand";
   attribute nokkelord of R50206 : Label is "Resistor Motstand";
   attribute nokkelord of R50205 : Label is "Resistor Motstand";
   attribute nokkelord of R50204 : Label is "Resistor Motstand";
   attribute nokkelord of R50203 : Label is "Resistor Motstand";
   attribute nokkelord of R50202 : Label is "Resistor Motstand";
   attribute nokkelord of R50201 : Label is "Resistor";
   attribute nokkelord of R50200 : Label is "Resistor";
   attribute nokkelord of J50206 : Label is "IDE";
   attribute nokkelord of J50205 : Label is "Connector, Kontakt";
   attribute nokkelord of J50204 : Label is "Connector, Kontakt";
   attribute nokkelord of J50203 : Label is "Connector, Kontakt";
   attribute nokkelord of J50202 : Label is "Connector, Kontakt";
   attribute nokkelord of J50201 : Label is "Connector, Kontakt";
   attribute nokkelord of J50200 : Label is "Connector, Kontakt";
   attribute nokkelord of D50217 : Label is "diode, led, lys, green";
   attribute nokkelord of D50215 : Label is "diode, led, lys, green";
   attribute nokkelord of D50214 : Label is "diode, led, lys, green";
   attribute nokkelord of D50212 : Label is "diode, led, lys, green";
   attribute nokkelord of D50211 : Label is "diode, led, lys, green";
   attribute nokkelord of D50209 : Label is "diode, led, lys, green";
   attribute nokkelord of D50208 : Label is "diode, led, lys, green";
   attribute nokkelord of D50206 : Label is "diode, led, lys, green";
   attribute nokkelord of D50205 : Label is "diode, led, lys, green";
   attribute nokkelord of D50203 : Label is "diode, led, lys, green";
   attribute nokkelord of D50202 : Label is "diode, led, lys, green";
   attribute nokkelord of D50200 : Label is "diode, led, lys, green";

   attribute pakke_opprettet : string;
   attribute pakke_opprettet of R50223 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50222 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50221 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50220 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50219 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50218 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50217 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50216 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50215 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50214 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50213 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50212 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50211 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50210 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50209 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50208 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50207 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50206 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50205 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50204 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50203 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50202 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50201 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of R50200 : Label is "08.07.2014 21:15:30";
   attribute pakke_opprettet of J50206 : Label is "12.07.2014 17.05.20";
   attribute pakke_opprettet of J50205 : Label is "28.06.2014 18:25:12";
   attribute pakke_opprettet of J50204 : Label is "28.06.2014 18:25:12";
   attribute pakke_opprettet of J50203 : Label is "28.06.2014 18:25:12";
   attribute pakke_opprettet of J50202 : Label is "28.06.2014 18:25:12";
   attribute pakke_opprettet of J50201 : Label is "28.06.2014 18:25:12";
   attribute pakke_opprettet of J50200 : Label is "28.06.2014 18:25:12";
   attribute pakke_opprettet of D50217 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50216 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50215 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50214 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50213 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50212 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50211 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50210 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50209 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50208 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50207 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50206 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50205 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50204 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50203 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50202 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50201 : Label is "09.02.2016 18:21:00";
   attribute pakke_opprettet of D50200 : Label is "09.02.2016 18:21:00";

   attribute pakke_opprettet_av : string;
   attribute pakke_opprettet_av of R50223 : Label is "815";
   attribute pakke_opprettet_av of R50222 : Label is "815";
   attribute pakke_opprettet_av of R50221 : Label is "815";
   attribute pakke_opprettet_av of R50220 : Label is "815";
   attribute pakke_opprettet_av of R50219 : Label is "815";
   attribute pakke_opprettet_av of R50218 : Label is "815";
   attribute pakke_opprettet_av of R50217 : Label is "815";
   attribute pakke_opprettet_av of R50216 : Label is "815";
   attribute pakke_opprettet_av of R50215 : Label is "815";
   attribute pakke_opprettet_av of R50214 : Label is "815";
   attribute pakke_opprettet_av of R50213 : Label is "815";
   attribute pakke_opprettet_av of R50212 : Label is "815";
   attribute pakke_opprettet_av of R50211 : Label is "815";
   attribute pakke_opprettet_av of R50210 : Label is "815";
   attribute pakke_opprettet_av of R50209 : Label is "815";
   attribute pakke_opprettet_av of R50208 : Label is "815";
   attribute pakke_opprettet_av of R50207 : Label is "815";
   attribute pakke_opprettet_av of R50206 : Label is "815";
   attribute pakke_opprettet_av of R50205 : Label is "815";
   attribute pakke_opprettet_av of R50204 : Label is "815";
   attribute pakke_opprettet_av of R50203 : Label is "815";
   attribute pakke_opprettet_av of R50202 : Label is "815";
   attribute pakke_opprettet_av of R50201 : Label is "815";
   attribute pakke_opprettet_av of R50200 : Label is "815";
   attribute pakke_opprettet_av of J50206 : Label is "815";
   attribute pakke_opprettet_av of J50205 : Label is "815";
   attribute pakke_opprettet_av of J50204 : Label is "815";
   attribute pakke_opprettet_av of J50203 : Label is "815";
   attribute pakke_opprettet_av of J50202 : Label is "815";
   attribute pakke_opprettet_av of J50201 : Label is "815";
   attribute pakke_opprettet_av of J50200 : Label is "815";
   attribute pakke_opprettet_av of D50217 : Label is "1366";
   attribute pakke_opprettet_av of D50216 : Label is "1366";
   attribute pakke_opprettet_av of D50215 : Label is "1366";
   attribute pakke_opprettet_av of D50214 : Label is "1366";
   attribute pakke_opprettet_av of D50213 : Label is "1366";
   attribute pakke_opprettet_av of D50212 : Label is "1366";
   attribute pakke_opprettet_av of D50211 : Label is "1366";
   attribute pakke_opprettet_av of D50210 : Label is "1366";
   attribute pakke_opprettet_av of D50209 : Label is "1366";
   attribute pakke_opprettet_av of D50208 : Label is "1366";
   attribute pakke_opprettet_av of D50207 : Label is "1366";
   attribute pakke_opprettet_av of D50206 : Label is "1366";
   attribute pakke_opprettet_av of D50205 : Label is "1366";
   attribute pakke_opprettet_av of D50204 : Label is "1366";
   attribute pakke_opprettet_av of D50203 : Label is "1366";
   attribute pakke_opprettet_av of D50202 : Label is "1366";
   attribute pakke_opprettet_av of D50201 : Label is "1366";
   attribute pakke_opprettet_av of D50200 : Label is "1366";

   attribute pakketype : string;
   attribute pakketype of R50223 : Label is "0603";
   attribute pakketype of R50222 : Label is "0603";
   attribute pakketype of R50221 : Label is "0603";
   attribute pakketype of R50220 : Label is "0603";
   attribute pakketype of R50219 : Label is "0603";
   attribute pakketype of R50218 : Label is "0603";
   attribute pakketype of R50217 : Label is "0603";
   attribute pakketype of R50216 : Label is "0603";
   attribute pakketype of R50215 : Label is "0603";
   attribute pakketype of R50214 : Label is "0603";
   attribute pakketype of R50213 : Label is "0603";
   attribute pakketype of R50212 : Label is "0603";
   attribute pakketype of R50211 : Label is "0603";
   attribute pakketype of R50210 : Label is "0603";
   attribute pakketype of R50209 : Label is "0603";
   attribute pakketype of R50208 : Label is "0603";
   attribute pakketype of R50207 : Label is "0603";
   attribute pakketype of R50206 : Label is "0603";
   attribute pakketype of R50205 : Label is "0603";
   attribute pakketype of R50204 : Label is "0603";
   attribute pakketype of R50203 : Label is "0603";
   attribute pakketype of R50202 : Label is "0603";
   attribute pakketype of R50201 : Label is "0603";
   attribute pakketype of R50200 : Label is "0603";
   attribute pakketype of J50206 : Label is "TH";
   attribute pakketype of J50205 : Label is "TH";
   attribute pakketype of J50204 : Label is "TH";
   attribute pakketype of J50203 : Label is "TH";
   attribute pakketype of J50202 : Label is "TH";
   attribute pakketype of J50201 : Label is "TH";
   attribute pakketype of J50200 : Label is "TH";
   attribute pakketype of D50217 : Label is "TH";
   attribute pakketype of D50216 : Label is "TH";
   attribute pakketype of D50215 : Label is "TH";
   attribute pakketype of D50214 : Label is "TH";
   attribute pakketype of D50213 : Label is "TH";
   attribute pakketype of D50212 : Label is "TH";
   attribute pakketype of D50211 : Label is "TH";
   attribute pakketype of D50210 : Label is "TH";
   attribute pakketype of D50209 : Label is "TH";
   attribute pakketype of D50208 : Label is "TH";
   attribute pakketype of D50207 : Label is "TH";
   attribute pakketype of D50206 : Label is "TH";
   attribute pakketype of D50205 : Label is "TH";
   attribute pakketype of D50204 : Label is "TH";
   attribute pakketype of D50203 : Label is "TH";
   attribute pakketype of D50202 : Label is "TH";
   attribute pakketype of D50201 : Label is "TH";
   attribute pakketype of D50200 : Label is "TH";

   attribute pris : string;
   attribute pris of R50223 : Label is "0";
   attribute pris of R50222 : Label is "0";
   attribute pris of R50221 : Label is "0";
   attribute pris of R50220 : Label is "0";
   attribute pris of R50219 : Label is "0";
   attribute pris of R50218 : Label is "0";
   attribute pris of R50217 : Label is "0";
   attribute pris of R50216 : Label is "0";
   attribute pris of R50215 : Label is "0";
   attribute pris of R50214 : Label is "0";
   attribute pris of R50213 : Label is "0";
   attribute pris of R50212 : Label is "0";
   attribute pris of R50211 : Label is "0";
   attribute pris of R50210 : Label is "0";
   attribute pris of R50209 : Label is "0";
   attribute pris of R50208 : Label is "0";
   attribute pris of R50207 : Label is "0";
   attribute pris of R50206 : Label is "0";
   attribute pris of R50205 : Label is "0";
   attribute pris of R50204 : Label is "0";
   attribute pris of R50203 : Label is "0";
   attribute pris of R50202 : Label is "0";
   attribute pris of R50201 : Label is "0";
   attribute pris of R50200 : Label is "0";
   attribute pris of J50206 : Label is "10";
   attribute pris of J50205 : Label is "2";
   attribute pris of J50204 : Label is "2";
   attribute pris of J50203 : Label is "2";
   attribute pris of J50202 : Label is "2";
   attribute pris of J50201 : Label is "2";
   attribute pris of J50200 : Label is "2";
   attribute pris of D50217 : Label is "3";
   attribute pris of D50216 : Label is "3";
   attribute pris of D50215 : Label is "3";
   attribute pris of D50214 : Label is "3";
   attribute pris of D50213 : Label is "3";
   attribute pris of D50212 : Label is "3";
   attribute pris of D50211 : Label is "3";
   attribute pris of D50210 : Label is "3";
   attribute pris of D50209 : Label is "3";
   attribute pris of D50208 : Label is "3";
   attribute pris of D50207 : Label is "3";
   attribute pris of D50206 : Label is "3";
   attribute pris of D50205 : Label is "3";
   attribute pris of D50204 : Label is "3";
   attribute pris of D50203 : Label is "3";
   attribute pris of D50202 : Label is "3";
   attribute pris of D50201 : Label is "3";
   attribute pris of D50200 : Label is "3";

   attribute produsent : string;
   attribute produsent of D50217 : Label is "Multikomp";
   attribute produsent of D50216 : Label is "Multicomp";
   attribute produsent of D50215 : Label is "Multikomp";
   attribute produsent of D50214 : Label is "Multikomp";
   attribute produsent of D50213 : Label is "Multicomp";
   attribute produsent of D50212 : Label is "Multikomp";
   attribute produsent of D50211 : Label is "Multikomp";
   attribute produsent of D50210 : Label is "Multicomp";
   attribute produsent of D50209 : Label is "Multikomp";
   attribute produsent of D50208 : Label is "Multikomp";
   attribute produsent of D50207 : Label is "Multicomp";
   attribute produsent of D50206 : Label is "Multikomp";
   attribute produsent of D50205 : Label is "Multikomp";
   attribute produsent of D50204 : Label is "Multicomp";
   attribute produsent of D50203 : Label is "Multikomp";
   attribute produsent of D50202 : Label is "Multikomp";
   attribute produsent of D50201 : Label is "Multicomp";
   attribute produsent of D50200 : Label is "Multikomp";

   attribute rad : string;
   attribute rad of R50223 : Label is "-1";
   attribute rad of R50222 : Label is "-1";
   attribute rad of R50221 : Label is "-1";
   attribute rad of R50220 : Label is "-1";
   attribute rad of R50219 : Label is "-1";
   attribute rad of R50218 : Label is "-1";
   attribute rad of R50217 : Label is "-1";
   attribute rad of R50216 : Label is "-1";
   attribute rad of R50215 : Label is "-1";
   attribute rad of R50214 : Label is "-1";
   attribute rad of R50213 : Label is "-1";
   attribute rad of R50212 : Label is "-1";
   attribute rad of R50211 : Label is "-1";
   attribute rad of R50210 : Label is "-1";
   attribute rad of R50209 : Label is "-1";
   attribute rad of R50208 : Label is "-1";
   attribute rad of R50207 : Label is "-1";
   attribute rad of R50206 : Label is "-1";
   attribute rad of R50205 : Label is "-1";
   attribute rad of R50204 : Label is "-1";
   attribute rad of R50203 : Label is "-1";
   attribute rad of R50202 : Label is "-1";
   attribute rad of R50201 : Label is "-1";
   attribute rad of R50200 : Label is "-1";

   attribute rom : string;
   attribute rom of R50223 : Label is "OV";
   attribute rom of R50222 : Label is "OV";
   attribute rom of R50221 : Label is "OV";
   attribute rom of R50220 : Label is "OV";
   attribute rom of R50219 : Label is "OV";
   attribute rom of R50218 : Label is "OV";
   attribute rom of R50217 : Label is "OV";
   attribute rom of R50216 : Label is "OV";
   attribute rom of R50215 : Label is "OV";
   attribute rom of R50214 : Label is "OV";
   attribute rom of R50213 : Label is "OV";
   attribute rom of R50212 : Label is "OV";
   attribute rom of R50211 : Label is "OV";
   attribute rom of R50210 : Label is "OV";
   attribute rom of R50209 : Label is "OV";
   attribute rom of R50208 : Label is "OV";
   attribute rom of R50207 : Label is "OV";
   attribute rom of R50206 : Label is "OV";
   attribute rom of R50205 : Label is "OV";
   attribute rom of R50204 : Label is "OV";
   attribute rom of R50203 : Label is "OV";
   attribute rom of R50202 : Label is "OV";
   attribute rom of R50201 : Label is "OV";
   attribute rom of R50200 : Label is "OV";

   attribute symbol_opprettet : string;
   attribute symbol_opprettet of R50223 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50222 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50221 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50220 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50219 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50218 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50217 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50216 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50215 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50214 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50213 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50212 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50211 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50210 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50209 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50208 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50207 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50206 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50205 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50204 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50203 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50202 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50201 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of R50200 : Label is "08.07.2014 21:16:33";
   attribute symbol_opprettet of J50206 : Label is "12.07.2014 17.03.56";
   attribute symbol_opprettet of J50205 : Label is "28.06.2014 15:33:24";
   attribute symbol_opprettet of J50204 : Label is "28.06.2014 15:33:24";
   attribute symbol_opprettet of J50203 : Label is "28.06.2014 15:33:24";
   attribute symbol_opprettet of J50202 : Label is "28.06.2014 15:33:24";
   attribute symbol_opprettet of J50201 : Label is "28.06.2014 15:33:24";
   attribute symbol_opprettet of J50200 : Label is "28.06.2014 15:33:24";
   attribute symbol_opprettet of D50217 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50216 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50215 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50214 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50213 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50212 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50211 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50210 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50209 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50208 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50207 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50206 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50205 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50204 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50203 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50202 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50201 : Label is "06.07.2014 18:59:47";
   attribute symbol_opprettet of D50200 : Label is "06.07.2014 18:59:47";

   attribute symbol_opprettet_av : string;
   attribute symbol_opprettet_av of R50223 : Label is "815";
   attribute symbol_opprettet_av of R50222 : Label is "815";
   attribute symbol_opprettet_av of R50221 : Label is "815";
   attribute symbol_opprettet_av of R50220 : Label is "815";
   attribute symbol_opprettet_av of R50219 : Label is "815";
   attribute symbol_opprettet_av of R50218 : Label is "815";
   attribute symbol_opprettet_av of R50217 : Label is "815";
   attribute symbol_opprettet_av of R50216 : Label is "815";
   attribute symbol_opprettet_av of R50215 : Label is "815";
   attribute symbol_opprettet_av of R50214 : Label is "815";
   attribute symbol_opprettet_av of R50213 : Label is "815";
   attribute symbol_opprettet_av of R50212 : Label is "815";
   attribute symbol_opprettet_av of R50211 : Label is "815";
   attribute symbol_opprettet_av of R50210 : Label is "815";
   attribute symbol_opprettet_av of R50209 : Label is "815";
   attribute symbol_opprettet_av of R50208 : Label is "815";
   attribute symbol_opprettet_av of R50207 : Label is "815";
   attribute symbol_opprettet_av of R50206 : Label is "815";
   attribute symbol_opprettet_av of R50205 : Label is "815";
   attribute symbol_opprettet_av of R50204 : Label is "815";
   attribute symbol_opprettet_av of R50203 : Label is "815";
   attribute symbol_opprettet_av of R50202 : Label is "815";
   attribute symbol_opprettet_av of R50201 : Label is "815";
   attribute symbol_opprettet_av of R50200 : Label is "815";
   attribute symbol_opprettet_av of J50206 : Label is "815";
   attribute symbol_opprettet_av of J50205 : Label is "815";
   attribute symbol_opprettet_av of J50204 : Label is "815";
   attribute symbol_opprettet_av of J50203 : Label is "815";
   attribute symbol_opprettet_av of J50202 : Label is "815";
   attribute symbol_opprettet_av of J50201 : Label is "815";
   attribute symbol_opprettet_av of J50200 : Label is "815";
   attribute symbol_opprettet_av of D50217 : Label is "815";
   attribute symbol_opprettet_av of D50216 : Label is "815";
   attribute symbol_opprettet_av of D50215 : Label is "815";
   attribute symbol_opprettet_av of D50214 : Label is "815";
   attribute symbol_opprettet_av of D50213 : Label is "815";
   attribute symbol_opprettet_av of D50212 : Label is "815";
   attribute symbol_opprettet_av of D50211 : Label is "815";
   attribute symbol_opprettet_av of D50210 : Label is "815";
   attribute symbol_opprettet_av of D50209 : Label is "815";
   attribute symbol_opprettet_av of D50208 : Label is "815";
   attribute symbol_opprettet_av of D50207 : Label is "815";
   attribute symbol_opprettet_av of D50206 : Label is "815";
   attribute symbol_opprettet_av of D50205 : Label is "815";
   attribute symbol_opprettet_av of D50204 : Label is "815";
   attribute symbol_opprettet_av of D50203 : Label is "815";
   attribute symbol_opprettet_av of D50202 : Label is "815";
   attribute symbol_opprettet_av of D50201 : Label is "815";
   attribute symbol_opprettet_av of D50200 : Label is "815";


Begin
    R50223 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50223|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50217_1,                           -- ObjectKind=Pin|PrimaryId=R50223-1
        X_2 => NamedSignal_5_ST                              -- ObjectKind=Pin|PrimaryId=R50223-2
      );

    R50222 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50222|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50216_1,                           -- ObjectKind=Pin|PrimaryId=R50222-1
        X_2 => NamedSignal_5_FE                              -- ObjectKind=Pin|PrimaryId=R50222-2
      );

    R50221 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50221|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50215_1,                           -- ObjectKind=Pin|PrimaryId=R50221-1
        X_2 => NamedSignal_5_KI                              -- ObjectKind=Pin|PrimaryId=R50221-2
      );

    R50220 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50220|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50214_1,                           -- ObjectKind=Pin|PrimaryId=R50220-1
        X_2 => NamedSignal_4_ST                              -- ObjectKind=Pin|PrimaryId=R50220-2
      );

    R50219 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50219|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50213_1,                           -- ObjectKind=Pin|PrimaryId=R50219-1
        X_2 => NamedSignal_4_FE                              -- ObjectKind=Pin|PrimaryId=R50219-2
      );

    R50218 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50218|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50212_1,                           -- ObjectKind=Pin|PrimaryId=R50218-1
        X_2 => NamedSignal_4_KI                              -- ObjectKind=Pin|PrimaryId=R50218-2
      );

    R50217 : X_2384                                          -- ObjectKind=Part|PrimaryId=R50217|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_5_KNP,                            -- ObjectKind=Pin|PrimaryId=R50217-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R50217-2
      );

    R50216 : X_2384                                          -- ObjectKind=Part|PrimaryId=R50216|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_4_KNP,                            -- ObjectKind=Pin|PrimaryId=R50216-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R50216-2
      );

    R50215 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50215|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50211_1,                           -- ObjectKind=Pin|PrimaryId=R50215-1
        X_2 => NamedSignal_3_ST                              -- ObjectKind=Pin|PrimaryId=R50215-2
      );

    R50214 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50214|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50210_1,                           -- ObjectKind=Pin|PrimaryId=R50214-1
        X_2 => NamedSignal_3_FE                              -- ObjectKind=Pin|PrimaryId=R50214-2
      );

    R50213 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50213|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50209_1,                           -- ObjectKind=Pin|PrimaryId=R50213-1
        X_2 => NamedSignal_3_KI                              -- ObjectKind=Pin|PrimaryId=R50213-2
      );

    R50212 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50212|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50208_1,                           -- ObjectKind=Pin|PrimaryId=R50212-1
        X_2 => NamedSignal_2_ST                              -- ObjectKind=Pin|PrimaryId=R50212-2
      );

    R50211 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50211|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50207_1,                           -- ObjectKind=Pin|PrimaryId=R50211-1
        X_2 => NamedSignal_2_FE                              -- ObjectKind=Pin|PrimaryId=R50211-2
      );

    R50210 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50210|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50206_1,                           -- ObjectKind=Pin|PrimaryId=R50210-1
        X_2 => NamedSignal_2_KI                              -- ObjectKind=Pin|PrimaryId=R50210-2
      );

    R50209 : X_2384                                          -- ObjectKind=Part|PrimaryId=R50209|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_3_KNP,                            -- ObjectKind=Pin|PrimaryId=R50209-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R50209-2
      );

    R50208 : X_2384                                          -- ObjectKind=Part|PrimaryId=R50208|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_2_KNP,                            -- ObjectKind=Pin|PrimaryId=R50208-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R50208-2
      );

    R50207 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50207|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50205_1,                           -- ObjectKind=Pin|PrimaryId=R50207-1
        X_2 => NamedSignal_1_ST                              -- ObjectKind=Pin|PrimaryId=R50207-2
      );

    R50206 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50206|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50204_1,                           -- ObjectKind=Pin|PrimaryId=R50206-1
        X_2 => NamedSignal_1_FE                              -- ObjectKind=Pin|PrimaryId=R50206-2
      );

    R50205 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50205|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50203_1,                           -- ObjectKind=Pin|PrimaryId=R50205-1
        X_2 => NamedSignal_1_KI                              -- ObjectKind=Pin|PrimaryId=R50205-2
      );

    R50204 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50204|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50202_1,                           -- ObjectKind=Pin|PrimaryId=R50204-1
        X_2 => NamedSignal_0_ST                              -- ObjectKind=Pin|PrimaryId=R50204-2
      );

    R50203 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50203|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50201_1,                           -- ObjectKind=Pin|PrimaryId=R50203-1
        X_2 => NamedSignal_0_FE                              -- ObjectKind=Pin|PrimaryId=R50203-2
      );

    R50202 : X_2448                                          -- ObjectKind=Part|PrimaryId=R50202|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50200_1,                           -- ObjectKind=Pin|PrimaryId=R50202-1
        X_2 => NamedSignal_0_KI                              -- ObjectKind=Pin|PrimaryId=R50202-2
      );

    R50201 : X_2384                                          -- ObjectKind=Part|PrimaryId=R50201|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_1_KNP,                            -- ObjectKind=Pin|PrimaryId=R50201-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R50201-2
      );

    R50200 : X_2384                                          -- ObjectKind=Part|PrimaryId=R50200|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_0_KNP,                            -- ObjectKind=Pin|PrimaryId=R50200-1
        X_2 => PowerSignal_VCC_P5V0                          -- ObjectKind=Pin|PrimaryId=R50200-2
      );

    J50206 : X_2390                                          -- ObjectKind=Part|PrimaryId=J50206|SecondaryId=1
      Port Map
      (
        X_1  => NamedSignal_0_KI,                            -- ObjectKind=Pin|PrimaryId=J50206-1
        X_2  => NamedSignal_1_KI,                            -- ObjectKind=Pin|PrimaryId=J50206-2
        X_3  => NamedSignal_0_FE,                            -- ObjectKind=Pin|PrimaryId=J50206-3
        X_4  => NamedSignal_1_FE,                            -- ObjectKind=Pin|PrimaryId=J50206-4
        X_5  => NamedSignal_0_ST,                            -- ObjectKind=Pin|PrimaryId=J50206-5
        X_6  => NamedSignal_1_ST,                            -- ObjectKind=Pin|PrimaryId=J50206-6
        X_7  => NamedSignal_0_INT,                           -- ObjectKind=Pin|PrimaryId=J50206-7
        X_8  => NamedSignal_1_INT,                           -- ObjectKind=Pin|PrimaryId=J50206-8
        X_9  => NamedSignal_0_KNP,                           -- ObjectKind=Pin|PrimaryId=J50206-9
        X_10 => NamedSignal_1_KNP,                           -- ObjectKind=Pin|PrimaryId=J50206-10
        X_11 => NamedSignal_2_KI,                            -- ObjectKind=Pin|PrimaryId=J50206-11
        X_12 => NamedSignal_3_KI,                            -- ObjectKind=Pin|PrimaryId=J50206-12
        X_13 => NamedSignal_2_FE,                            -- ObjectKind=Pin|PrimaryId=J50206-13
        X_14 => NamedSignal_3_FE,                            -- ObjectKind=Pin|PrimaryId=J50206-14
        X_15 => NamedSignal_2_ST,                            -- ObjectKind=Pin|PrimaryId=J50206-15
        X_16 => NamedSignal_3_ST,                            -- ObjectKind=Pin|PrimaryId=J50206-16
        X_17 => NamedSignal_2_INT,                           -- ObjectKind=Pin|PrimaryId=J50206-17
        X_18 => NamedSignal_3_INT,                           -- ObjectKind=Pin|PrimaryId=J50206-18
        X_19 => NamedSignal_2_KNP,                           -- ObjectKind=Pin|PrimaryId=J50206-19
        X_20 => NamedSignal_3_KNP,                           -- ObjectKind=Pin|PrimaryId=J50206-20
        X_21 => NamedSignal_4_KI,                            -- ObjectKind=Pin|PrimaryId=J50206-21
        X_22 => NamedSignal_5_KI,                            -- ObjectKind=Pin|PrimaryId=J50206-22
        X_23 => NamedSignal_4_FE,                            -- ObjectKind=Pin|PrimaryId=J50206-23
        X_24 => NamedSignal_5_FE,                            -- ObjectKind=Pin|PrimaryId=J50206-24
        X_25 => NamedSignal_4_ST,                            -- ObjectKind=Pin|PrimaryId=J50206-25
        X_26 => NamedSignal_5_ST,                            -- ObjectKind=Pin|PrimaryId=J50206-26
        X_27 => NamedSignal_4_INT,                           -- ObjectKind=Pin|PrimaryId=J50206-27
        X_28 => NamedSignal_5_INT,                           -- ObjectKind=Pin|PrimaryId=J50206-28
        X_29 => NamedSignal_4_KNP,                           -- ObjectKind=Pin|PrimaryId=J50206-29
        X_30 => NamedSignal_5_KNP,                           -- ObjectKind=Pin|PrimaryId=J50206-30
        X_31 => PowerSignal_VCC_P5V0,                        -- ObjectKind=Pin|PrimaryId=J50206-31
        X_32 => PowerSignal_GND,                             -- ObjectKind=Pin|PrimaryId=J50206-32
        X_33 => PowerSignal_VCC_P5V0,                        -- ObjectKind=Pin|PrimaryId=J50206-33
        X_34 => PowerSignal_GND                              -- ObjectKind=Pin|PrimaryId=J50206-34
      );

    J50205 : X_2226                                          -- ObjectKind=Part|PrimaryId=J50205|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_5_INT,                            -- ObjectKind=Pin|PrimaryId=J50205-1
        X_2 => NamedSignal_5_KNP,                            -- ObjectKind=Pin|PrimaryId=J50205-2
        X_3 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J50205-3
      );

    J50204 : X_2226                                          -- ObjectKind=Part|PrimaryId=J50204|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_4_INT,                            -- ObjectKind=Pin|PrimaryId=J50204-1
        X_2 => NamedSignal_4_KNP,                            -- ObjectKind=Pin|PrimaryId=J50204-2
        X_3 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J50204-3
      );

    J50203 : X_2226                                          -- ObjectKind=Part|PrimaryId=J50203|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_3_INT,                            -- ObjectKind=Pin|PrimaryId=J50203-1
        X_2 => NamedSignal_3_KNP,                            -- ObjectKind=Pin|PrimaryId=J50203-2
        X_3 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J50203-3
      );

    J50202 : X_2226                                          -- ObjectKind=Part|PrimaryId=J50202|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_2_INT,                            -- ObjectKind=Pin|PrimaryId=J50202-1
        X_2 => NamedSignal_2_KNP,                            -- ObjectKind=Pin|PrimaryId=J50202-2
        X_3 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J50202-3
      );

    J50201 : X_2226                                          -- ObjectKind=Part|PrimaryId=J50201|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_1_INT,                            -- ObjectKind=Pin|PrimaryId=J50201-1
        X_2 => NamedSignal_1_KNP,                            -- ObjectKind=Pin|PrimaryId=J50201-2
        X_3 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J50201-3
      );

    J50200 : X_2226                                          -- ObjectKind=Part|PrimaryId=J50200|SecondaryId=1
      Port Map
      (
        X_1 => NamedSignal_0_INT,                            -- ObjectKind=Pin|PrimaryId=J50200-1
        X_2 => NamedSignal_0_KNP,                            -- ObjectKind=Pin|PrimaryId=J50200-2
        X_3 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=J50200-3
      );

    D50217 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50217|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50217_1,                           -- ObjectKind=Pin|PrimaryId=D50217-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50217-2
      );

    D50216 : X_3597                                          -- ObjectKind=Part|PrimaryId=D50216|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50216_1,                           -- ObjectKind=Pin|PrimaryId=D50216-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50216-2
      );

    D50215 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50215|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50215_1,                           -- ObjectKind=Pin|PrimaryId=D50215-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50215-2
      );

    D50214 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50214|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50214_1,                           -- ObjectKind=Pin|PrimaryId=D50214-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50214-2
      );

    D50213 : X_3597                                          -- ObjectKind=Part|PrimaryId=D50213|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50213_1,                           -- ObjectKind=Pin|PrimaryId=D50213-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50213-2
      );

    D50212 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50212|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50212_1,                           -- ObjectKind=Pin|PrimaryId=D50212-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50212-2
      );

    D50211 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50211|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50211_1,                           -- ObjectKind=Pin|PrimaryId=D50211-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50211-2
      );

    D50210 : X_3597                                          -- ObjectKind=Part|PrimaryId=D50210|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50210_1,                           -- ObjectKind=Pin|PrimaryId=D50210-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50210-2
      );

    D50209 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50209|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50209_1,                           -- ObjectKind=Pin|PrimaryId=D50209-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50209-2
      );

    D50208 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50208|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50208_1,                           -- ObjectKind=Pin|PrimaryId=D50208-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50208-2
      );

    D50207 : X_3597                                          -- ObjectKind=Part|PrimaryId=D50207|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50207_1,                           -- ObjectKind=Pin|PrimaryId=D50207-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50207-2
      );

    D50206 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50206|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50206_1,                           -- ObjectKind=Pin|PrimaryId=D50206-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50206-2
      );

    D50205 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50205|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50205_1,                           -- ObjectKind=Pin|PrimaryId=D50205-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50205-2
      );

    D50204 : X_3597                                          -- ObjectKind=Part|PrimaryId=D50204|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50204_1,                           -- ObjectKind=Pin|PrimaryId=D50204-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50204-2
      );

    D50203 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50203|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50203_1,                           -- ObjectKind=Pin|PrimaryId=D50203-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50203-2
      );

    D50202 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50202|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50202_1,                           -- ObjectKind=Pin|PrimaryId=D50202-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50202-2
      );

    D50201 : X_3597                                          -- ObjectKind=Part|PrimaryId=D50201|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50201_1,                           -- ObjectKind=Pin|PrimaryId=D50201-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50201-2
      );

    D50200 : X_2076                                          -- ObjectKind=Part|PrimaryId=D50200|SecondaryId=1
      Port Map
      (
        X_1 => PinSignal_D50200_1,                           -- ObjectKind=Pin|PrimaryId=D50200-1
        X_2 => PowerSignal_GND                               -- ObjectKind=Pin|PrimaryId=D50200-2
      );

    -- Signal Assignments
    ---------------------
    PowerSignal_GND <= '0'; -- ObjectKind=Net|PrimaryId=GND

End Structure;
------------------------------------------------------------

