------------------------------------------------------------
-- VHDL TK532_Utgangskondensator
-- 2015 7 5 14 55 24
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 15.0.7.36915
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK532_Utgangskondensator
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK532_Utgangskondensator Is
  attribute MacroCell : boolean;

End TK532_Utgangskondensator;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK532_Utgangskondensator Is


Begin
End Structure;
------------------------------------------------------------

