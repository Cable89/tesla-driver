------------------------------------------------------------
-- VHDL TK516_EKSTRAMINUSPSU
-- 2014 7 8 19 13 37
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK516_EKSTRAMINUSPSU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK516_EKSTRAMINUSPSU Is
  attribute MacroCell : boolean;

End TK516_EKSTRAMINUSPSU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK516_EKSTRAMINUSPSU Is


Begin
End Structure;
------------------------------------------------------------

