------------------------------------------------------------
-- VHDL TK518_P18VMINUSPSU
-- 2017 1 13 17 4 7
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.0.6.282
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK518_P18VMINUSPSU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK518_P18VMINUSPSU Is
  attribute MacroCell : boolean;

End TK518_P18VMINUSPSU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK518_P18VMINUSPSU Is


Begin
End Structure;
------------------------------------------------------------

