------------------------------------------------------------
-- VHDL TK510_Mekanisk
-- 2014 7 12 21 47 5
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK510_Mekanisk
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK510_Mekanisk Is
  attribute MacroCell : boolean;

End TK510_Mekanisk;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK510_Mekanisk Is
   Component KortSt_tte                                      -- ObjectKind=Part|PrimaryId=M1|SecondaryId=1
   End Component;



   attribute antall : string;
   attribute antall of M18 : Label is "30";
   attribute antall of M17 : Label is "30";
   attribute antall of M16 : Label is "30";
   attribute antall of M15 : Label is "30";
   attribute antall of M14 : Label is "30";
   attribute antall of M13 : Label is "30";
   attribute antall of M12 : Label is "30";
   attribute antall of M11 : Label is "30";
   attribute antall of M10 : Label is "30";
   attribute antall of M9  : Label is "30";
   attribute antall of M8  : Label is "30";
   attribute antall of M7  : Label is "30";
   attribute antall of M6  : Label is "30";
   attribute antall of M5  : Label is "30";
   attribute antall of M4  : Label is "30";
   attribute antall of M3  : Label is "30";
   attribute antall of M2  : Label is "30";
   attribute antall of M1  : Label is "30";

   attribute beskrivelse : string;
   attribute beskrivelse of M18 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M17 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M16 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M15 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M14 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M13 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M12 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M11 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M10 : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M9  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M8  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M7  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M6  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M5  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M4  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M3  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M2  : Label is "St�tter kort i bakplan";
   attribute beskrivelse of M1  : Label is "St�tter kort i bakplan";

   attribute Database_Table_Name : string;
   attribute Database_Table_Name of M18 : Label is "altium";
   attribute Database_Table_Name of M17 : Label is "altium";
   attribute Database_Table_Name of M16 : Label is "altium";
   attribute Database_Table_Name of M15 : Label is "altium";
   attribute Database_Table_Name of M14 : Label is "altium";
   attribute Database_Table_Name of M13 : Label is "altium";
   attribute Database_Table_Name of M12 : Label is "altium";
   attribute Database_Table_Name of M11 : Label is "altium";
   attribute Database_Table_Name of M10 : Label is "altium";
   attribute Database_Table_Name of M9  : Label is "altium";
   attribute Database_Table_Name of M8  : Label is "altium";
   attribute Database_Table_Name of M7  : Label is "altium";
   attribute Database_Table_Name of M6  : Label is "altium";
   attribute Database_Table_Name of M5  : Label is "altium";
   attribute Database_Table_Name of M4  : Label is "altium";
   attribute Database_Table_Name of M3  : Label is "altium";
   attribute Database_Table_Name of M2  : Label is "altium";
   attribute Database_Table_Name of M1  : Label is "altium";

   attribute dybde : string;
   attribute dybde of M18 : Label is "0";
   attribute dybde of M17 : Label is "0";
   attribute dybde of M16 : Label is "0";
   attribute dybde of M15 : Label is "0";
   attribute dybde of M14 : Label is "0";
   attribute dybde of M13 : Label is "0";
   attribute dybde of M12 : Label is "0";
   attribute dybde of M11 : Label is "0";
   attribute dybde of M10 : Label is "0";
   attribute dybde of M9  : Label is "0";
   attribute dybde of M8  : Label is "0";
   attribute dybde of M7  : Label is "0";
   attribute dybde of M6  : Label is "0";
   attribute dybde of M5  : Label is "0";
   attribute dybde of M4  : Label is "0";
   attribute dybde of M3  : Label is "0";
   attribute dybde of M2  : Label is "0";
   attribute dybde of M1  : Label is "0";

   attribute hylle : string;
   attribute hylle of M18 : Label is "15";
   attribute hylle of M17 : Label is "15";
   attribute hylle of M16 : Label is "15";
   attribute hylle of M15 : Label is "15";
   attribute hylle of M14 : Label is "15";
   attribute hylle of M13 : Label is "15";
   attribute hylle of M12 : Label is "15";
   attribute hylle of M11 : Label is "15";
   attribute hylle of M10 : Label is "15";
   attribute hylle of M9  : Label is "15";
   attribute hylle of M8  : Label is "15";
   attribute hylle of M7  : Label is "15";
   attribute hylle of M6  : Label is "15";
   attribute hylle of M5  : Label is "15";
   attribute hylle of M4  : Label is "15";
   attribute hylle of M3  : Label is "15";
   attribute hylle of M2  : Label is "15";
   attribute hylle of M1  : Label is "15";

   attribute kolonne : string;
   attribute kolonne of M18 : Label is "2";
   attribute kolonne of M17 : Label is "2";
   attribute kolonne of M16 : Label is "2";
   attribute kolonne of M15 : Label is "2";
   attribute kolonne of M14 : Label is "2";
   attribute kolonne of M13 : Label is "2";
   attribute kolonne of M12 : Label is "2";
   attribute kolonne of M11 : Label is "2";
   attribute kolonne of M10 : Label is "2";
   attribute kolonne of M9  : Label is "2";
   attribute kolonne of M8  : Label is "2";
   attribute kolonne of M7  : Label is "2";
   attribute kolonne of M6  : Label is "2";
   attribute kolonne of M5  : Label is "2";
   attribute kolonne of M4  : Label is "2";
   attribute kolonne of M3  : Label is "2";
   attribute kolonne of M2  : Label is "2";
   attribute kolonne of M1  : Label is "2";

   attribute lager_type : string;
   attribute lager_type of M18 : Label is "Fremlager";
   attribute lager_type of M17 : Label is "Fremlager";
   attribute lager_type of M16 : Label is "Fremlager";
   attribute lager_type of M15 : Label is "Fremlager";
   attribute lager_type of M14 : Label is "Fremlager";
   attribute lager_type of M13 : Label is "Fremlager";
   attribute lager_type of M12 : Label is "Fremlager";
   attribute lager_type of M11 : Label is "Fremlager";
   attribute lager_type of M10 : Label is "Fremlager";
   attribute lager_type of M9  : Label is "Fremlager";
   attribute lager_type of M8  : Label is "Fremlager";
   attribute lager_type of M7  : Label is "Fremlager";
   attribute lager_type of M6  : Label is "Fremlager";
   attribute lager_type of M5  : Label is "Fremlager";
   attribute lager_type of M4  : Label is "Fremlager";
   attribute lager_type of M3  : Label is "Fremlager";
   attribute lager_type of M2  : Label is "Fremlager";
   attribute lager_type of M1  : Label is "Fremlager";

   attribute navn : string;
   attribute navn of M18 : Label is "KortSt�tte";
   attribute navn of M17 : Label is "KortSt�tte";
   attribute navn of M16 : Label is "KortSt�tte";
   attribute navn of M15 : Label is "KortSt�tte";
   attribute navn of M14 : Label is "KortSt�tte";
   attribute navn of M13 : Label is "KortSt�tte";
   attribute navn of M12 : Label is "KortSt�tte";
   attribute navn of M11 : Label is "KortSt�tte";
   attribute navn of M10 : Label is "KortSt�tte";
   attribute navn of M9  : Label is "KortSt�tte";
   attribute navn of M8  : Label is "KortSt�tte";
   attribute navn of M7  : Label is "KortSt�tte";
   attribute navn of M6  : Label is "KortSt�tte";
   attribute navn of M5  : Label is "KortSt�tte";
   attribute navn of M4  : Label is "KortSt�tte";
   attribute navn of M3  : Label is "KortSt�tte";
   attribute navn of M2  : Label is "KortSt�tte";
   attribute navn of M1  : Label is "KortSt�tte";

   attribute nokkelord : string;
   attribute nokkelord of M18 : Label is "support";
   attribute nokkelord of M17 : Label is "support";
   attribute nokkelord of M16 : Label is "support";
   attribute nokkelord of M15 : Label is "support";
   attribute nokkelord of M14 : Label is "support";
   attribute nokkelord of M13 : Label is "support";
   attribute nokkelord of M12 : Label is "support";
   attribute nokkelord of M11 : Label is "support";
   attribute nokkelord of M10 : Label is "support";
   attribute nokkelord of M9  : Label is "support";
   attribute nokkelord of M8  : Label is "support";
   attribute nokkelord of M7  : Label is "support";
   attribute nokkelord of M6  : Label is "support";
   attribute nokkelord of M5  : Label is "support";
   attribute nokkelord of M4  : Label is "support";
   attribute nokkelord of M3  : Label is "support";
   attribute nokkelord of M2  : Label is "support";
   attribute nokkelord of M1  : Label is "support";

   attribute pakke_opprettet : string;
   attribute pakke_opprettet of M18 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M17 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M16 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M15 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M14 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M13 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M12 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M11 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M10 : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M9  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M8  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M7  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M6  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M5  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M4  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M3  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M2  : Label is "12.07.2014 20:29:43";
   attribute pakke_opprettet of M1  : Label is "12.07.2014 20:29:43";

   attribute pakke_opprettet_av : string;
   attribute pakke_opprettet_av of M18 : Label is "815";
   attribute pakke_opprettet_av of M17 : Label is "815";
   attribute pakke_opprettet_av of M16 : Label is "815";
   attribute pakke_opprettet_av of M15 : Label is "815";
   attribute pakke_opprettet_av of M14 : Label is "815";
   attribute pakke_opprettet_av of M13 : Label is "815";
   attribute pakke_opprettet_av of M12 : Label is "815";
   attribute pakke_opprettet_av of M11 : Label is "815";
   attribute pakke_opprettet_av of M10 : Label is "815";
   attribute pakke_opprettet_av of M9  : Label is "815";
   attribute pakke_opprettet_av of M8  : Label is "815";
   attribute pakke_opprettet_av of M7  : Label is "815";
   attribute pakke_opprettet_av of M6  : Label is "815";
   attribute pakke_opprettet_av of M5  : Label is "815";
   attribute pakke_opprettet_av of M4  : Label is "815";
   attribute pakke_opprettet_av of M3  : Label is "815";
   attribute pakke_opprettet_av of M2  : Label is "815";
   attribute pakke_opprettet_av of M1  : Label is "815";

   attribute pakketype : string;
   attribute pakketype of M18 : Label is "92";
   attribute pakketype of M17 : Label is "92";
   attribute pakketype of M16 : Label is "92";
   attribute pakketype of M15 : Label is "92";
   attribute pakketype of M14 : Label is "92";
   attribute pakketype of M13 : Label is "92";
   attribute pakketype of M12 : Label is "92";
   attribute pakketype of M11 : Label is "92";
   attribute pakketype of M10 : Label is "92";
   attribute pakketype of M9  : Label is "92";
   attribute pakketype of M8  : Label is "92";
   attribute pakketype of M7  : Label is "92";
   attribute pakketype of M6  : Label is "92";
   attribute pakketype of M5  : Label is "92";
   attribute pakketype of M4  : Label is "92";
   attribute pakketype of M3  : Label is "92";
   attribute pakketype of M2  : Label is "92";
   attribute pakketype of M1  : Label is "92";

   attribute pris : string;
   attribute pris of M18 : Label is "5";
   attribute pris of M17 : Label is "5";
   attribute pris of M16 : Label is "5";
   attribute pris of M15 : Label is "5";
   attribute pris of M14 : Label is "5";
   attribute pris of M13 : Label is "5";
   attribute pris of M12 : Label is "5";
   attribute pris of M11 : Label is "5";
   attribute pris of M10 : Label is "5";
   attribute pris of M9  : Label is "5";
   attribute pris of M8  : Label is "5";
   attribute pris of M7  : Label is "5";
   attribute pris of M6  : Label is "5";
   attribute pris of M5  : Label is "5";
   attribute pris of M4  : Label is "5";
   attribute pris of M3  : Label is "5";
   attribute pris of M2  : Label is "5";
   attribute pris of M1  : Label is "5";

   attribute rad : string;
   attribute rad of M18 : Label is "5";
   attribute rad of M17 : Label is "5";
   attribute rad of M16 : Label is "5";
   attribute rad of M15 : Label is "5";
   attribute rad of M14 : Label is "5";
   attribute rad of M13 : Label is "5";
   attribute rad of M12 : Label is "5";
   attribute rad of M11 : Label is "5";
   attribute rad of M10 : Label is "5";
   attribute rad of M9  : Label is "5";
   attribute rad of M8  : Label is "5";
   attribute rad of M7  : Label is "5";
   attribute rad of M6  : Label is "5";
   attribute rad of M5  : Label is "5";
   attribute rad of M4  : Label is "5";
   attribute rad of M3  : Label is "5";
   attribute rad of M2  : Label is "5";
   attribute rad of M1  : Label is "5";

   attribute rom : string;
   attribute rom of M18 : Label is "OV";
   attribute rom of M17 : Label is "OV";
   attribute rom of M16 : Label is "OV";
   attribute rom of M15 : Label is "OV";
   attribute rom of M14 : Label is "OV";
   attribute rom of M13 : Label is "OV";
   attribute rom of M12 : Label is "OV";
   attribute rom of M11 : Label is "OV";
   attribute rom of M10 : Label is "OV";
   attribute rom of M9  : Label is "OV";
   attribute rom of M8  : Label is "OV";
   attribute rom of M7  : Label is "OV";
   attribute rom of M6  : Label is "OV";
   attribute rom of M5  : Label is "OV";
   attribute rom of M4  : Label is "OV";
   attribute rom of M3  : Label is "OV";
   attribute rom of M2  : Label is "OV";
   attribute rom of M1  : Label is "OV";

   attribute symbol_opprettet : string;
   attribute symbol_opprettet of M18 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M17 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M16 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M15 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M14 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M13 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M12 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M11 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M10 : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M9  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M8  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M7  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M6  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M5  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M4  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M3  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M2  : Label is "12.07.2014 20:29:53";
   attribute symbol_opprettet of M1  : Label is "12.07.2014 20:29:53";

   attribute symbol_opprettet_av : string;
   attribute symbol_opprettet_av of M18 : Label is "815";
   attribute symbol_opprettet_av of M17 : Label is "815";
   attribute symbol_opprettet_av of M16 : Label is "815";
   attribute symbol_opprettet_av of M15 : Label is "815";
   attribute symbol_opprettet_av of M14 : Label is "815";
   attribute symbol_opprettet_av of M13 : Label is "815";
   attribute symbol_opprettet_av of M12 : Label is "815";
   attribute symbol_opprettet_av of M11 : Label is "815";
   attribute symbol_opprettet_av of M10 : Label is "815";
   attribute symbol_opprettet_av of M9  : Label is "815";
   attribute symbol_opprettet_av of M8  : Label is "815";
   attribute symbol_opprettet_av of M7  : Label is "815";
   attribute symbol_opprettet_av of M6  : Label is "815";
   attribute symbol_opprettet_av of M5  : Label is "815";
   attribute symbol_opprettet_av of M4  : Label is "815";
   attribute symbol_opprettet_av of M3  : Label is "815";
   attribute symbol_opprettet_av of M2  : Label is "815";
   attribute symbol_opprettet_av of M1  : Label is "815";


Begin
    M18 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M18|SecondaryId=1
;

    M17 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M17|SecondaryId=1
;

    M16 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M16|SecondaryId=1
;

    M15 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M15|SecondaryId=1
;

    M14 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M14|SecondaryId=1
;

    M13 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M13|SecondaryId=1
;

    M12 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M12|SecondaryId=1
;

    M11 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M11|SecondaryId=1
;

    M10 : KortSt_tte                                         -- ObjectKind=Part|PrimaryId=M10|SecondaryId=1
;

    M9 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M9|SecondaryId=1
;

    M8 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M8|SecondaryId=1
;

    M7 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M7|SecondaryId=1
;

    M6 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M6|SecondaryId=1
;

    M5 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M5|SecondaryId=1
;

    M4 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M4|SecondaryId=1
;

    M3 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M3|SecondaryId=1
;

    M2 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M2|SecondaryId=1
;

    M1 : KortSt_tte                                          -- ObjectKind=Part|PrimaryId=M1|SecondaryId=1
;

End Structure;
------------------------------------------------------------

