------------------------------------------------------------
-- VHDL TK518_P18VMINUSPSU
-- 2014 7 12 21 38 42
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK518_P18VMINUSPSU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK518_P18VMINUSPSU Is
  attribute MacroCell : boolean;

End TK518_P18VMINUSPSU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK518_P18VMINUSPSU Is


Begin
End Structure;
------------------------------------------------------------

