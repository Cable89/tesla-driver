------------------------------------------------------------
-- VHDL TK511_Blindkort
-- 2014 7 12 21 38 42
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK511_Blindkort
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK511_Blindkort Is
  port
  (
    A1           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A1
    A2           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A2
    A3           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A3
    A4           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A4
    A5           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A5
    A6           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A6
    A7           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A7
    A8           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A8
    A9           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=A9
    B3           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B3
    B4           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B4
    B5           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B5
    B6           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B6
    B7           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B7
    B8           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B8
    B9           : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B9
    B10          : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B10
    B11          : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B11
    B12          : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B12
    B13          : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B13
    B14          : InOut STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=B14
    FEIL         : Out   STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=FEIL
    INTERRUPT    : Out   STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=INTERRUPT
    KORT_INNSATT : Out   STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=KORT INNSATT
    LIMIT        : In    STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=LIMIT
    RESERVELED   : Out   STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=RESERVELED
    STATUS       : Out   STD_LOGIC;                          -- ObjectKind=Port|PrimaryId=STATUS
    TRIGGER      : In    STD_LOGIC                           -- ObjectKind=Port|PrimaryId=TRIGGER
  );
  attribute MacroCell : boolean;

End TK511_Blindkort;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK511_Blindkort Is


Begin
End Structure;
------------------------------------------------------------

