------------------------------------------------------------
-- VHDL TK540_Frontpanel
-- 2014 7 8 19 13 37
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL TK540_Frontpanel
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity TK540_Frontpanel Is
  attribute MacroCell : boolean;

End TK540_Frontpanel;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of TK540_Frontpanel Is


Begin
End Structure;
------------------------------------------------------------

